* SPICE NETLIST
***************************************

.SUBCKT M1_POLY_CDNS_712283338712
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NTAP_CDNS_712283338711
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT PTAP_CDNS_712283338710
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_1
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_2
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_3
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_4
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_5
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_6
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_7
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_8
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_9
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_10
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_11
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_12
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_13
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_14
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_15
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_16
** N=1 EP=0 IP=3 FDC=0
.ENDS
***************************************
.SUBCKT ICV_17
** N=1 EP=0 IP=3 FDC=0
.ENDS
***************************************
.SUBCKT ICV_18
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_19
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_20
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_21
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_22
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_23
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_24 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165
** N=1091 EP=165 IP=2241 FDC=2700
M0 166 1 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=134870 $D=1
M1 167 1 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=139500 $D=1
M2 168 1 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=144130 $D=1
M3 169 166 2 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=134870 $D=1
M4 170 167 3 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=139500 $D=1
M5 171 168 4 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=144130 $D=1
M6 9 1 169 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=134870 $D=1
M7 9 1 170 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=139500 $D=1
M8 9 1 171 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=144130 $D=1
M9 172 166 2 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=134870 $D=1
M10 173 167 3 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=139500 $D=1
M11 174 168 4 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=144130 $D=1
M12 2 1 172 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=134870 $D=1
M13 3 1 173 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=139500 $D=1
M14 4 1 174 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=144130 $D=1
M15 175 166 2 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=134870 $D=1
M16 176 167 3 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=139500 $D=1
M17 177 168 4 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=144130 $D=1
M18 2 1 175 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=134870 $D=1
M19 3 1 176 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=139500 $D=1
M20 4 1 177 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=144130 $D=1
M21 181 178 175 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=134870 $D=1
M22 182 179 176 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=139500 $D=1
M23 183 180 177 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=144130 $D=1
M24 178 5 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=134870 $D=1
M25 179 5 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=139500 $D=1
M26 180 5 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=144130 $D=1
M27 184 178 172 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=134870 $D=1
M28 185 179 173 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=139500 $D=1
M29 186 180 174 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=144130 $D=1
M30 169 5 184 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=134870 $D=1
M31 170 5 185 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=139500 $D=1
M32 171 5 186 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=144130 $D=1
M33 187 6 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=134870 $D=1
M34 188 6 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=139500 $D=1
M35 189 6 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=144130 $D=1
M36 190 187 184 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=134870 $D=1
M37 191 188 185 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=139500 $D=1
M38 192 189 186 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=144130 $D=1
M39 181 6 190 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=134870 $D=1
M40 182 6 191 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=139500 $D=1
M41 183 6 192 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=144130 $D=1
M42 193 8 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=134870 $D=1
M43 194 8 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=139500 $D=1
M44 195 8 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=144130 $D=1
M45 196 193 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=134870 $D=1
M46 197 194 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=139500 $D=1
M47 198 195 10 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=144130 $D=1
M48 11 8 196 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=134870 $D=1
M49 12 8 197 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=139500 $D=1
M50 13 8 198 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=144130 $D=1
M51 199 193 14 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=134870 $D=1
M52 200 194 15 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=139500 $D=1
M53 201 195 16 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=144130 $D=1
M54 202 8 199 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=134870 $D=1
M55 203 8 200 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=139500 $D=1
M56 204 8 201 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=144130 $D=1
M57 208 193 205 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=134870 $D=1
M58 209 194 206 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=139500 $D=1
M59 210 195 207 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=144130 $D=1
M60 190 8 208 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=134870 $D=1
M61 191 8 209 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=139500 $D=1
M62 192 8 210 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=144130 $D=1
M63 214 211 208 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=134870 $D=1
M64 215 212 209 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=139500 $D=1
M65 216 213 210 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=144130 $D=1
M66 211 17 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=134870 $D=1
M67 212 17 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=139500 $D=1
M68 213 17 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=144130 $D=1
M69 217 211 199 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=134870 $D=1
M70 218 212 200 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=139500 $D=1
M71 219 213 201 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=144130 $D=1
M72 196 17 217 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=134870 $D=1
M73 197 17 218 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=139500 $D=1
M74 198 17 219 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=144130 $D=1
M75 220 18 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=134870 $D=1
M76 221 18 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=139500 $D=1
M77 222 18 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=144130 $D=1
M78 223 220 217 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=134870 $D=1
M79 224 221 218 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=139500 $D=1
M80 225 222 219 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=144130 $D=1
M81 214 18 223 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=134870 $D=1
M82 215 18 224 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=139500 $D=1
M83 216 18 225 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=144130 $D=1
M84 9 19 226 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=134870 $D=1
M85 9 19 227 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=139500 $D=1
M86 9 19 228 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=144130 $D=1
M87 229 20 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=134870 $D=1
M88 230 20 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=139500 $D=1
M89 231 20 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=144130 $D=1
M90 232 19 223 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=134870 $D=1
M91 233 19 224 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=139500 $D=1
M92 234 19 225 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=144130 $D=1
M93 9 232 939 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=134870 $D=1
M94 9 233 940 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=139500 $D=1
M95 9 234 941 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=144130 $D=1
M96 235 939 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=134870 $D=1
M97 236 940 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=139500 $D=1
M98 237 941 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=144130 $D=1
M99 232 226 235 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=134870 $D=1
M100 233 227 236 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=139500 $D=1
M101 234 228 237 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=144130 $D=1
M102 235 20 238 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=134870 $D=1
M103 236 20 239 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=139500 $D=1
M104 237 20 240 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=144130 $D=1
M105 244 21 235 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=134870 $D=1
M106 245 21 236 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=139500 $D=1
M107 246 21 237 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=144130 $D=1
M108 241 21 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=134870 $D=1
M109 242 21 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=139500 $D=1
M110 243 21 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=144130 $D=1
M111 9 22 247 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=134870 $D=1
M112 9 22 248 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=139500 $D=1
M113 9 22 249 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=144130 $D=1
M114 250 23 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=134870 $D=1
M115 251 23 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=139500 $D=1
M116 252 23 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=144130 $D=1
M117 253 22 223 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=134870 $D=1
M118 254 22 224 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=139500 $D=1
M119 255 22 225 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=144130 $D=1
M120 9 253 942 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=134870 $D=1
M121 9 254 943 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=139500 $D=1
M122 9 255 944 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=144130 $D=1
M123 256 942 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=134870 $D=1
M124 257 943 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=139500 $D=1
M125 258 944 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=144130 $D=1
M126 253 247 256 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=134870 $D=1
M127 254 248 257 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=139500 $D=1
M128 255 249 258 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=144130 $D=1
M129 256 23 238 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=134870 $D=1
M130 257 23 239 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=139500 $D=1
M131 258 23 240 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=144130 $D=1
M132 244 24 256 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=134870 $D=1
M133 245 24 257 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=139500 $D=1
M134 246 24 258 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=144130 $D=1
M135 259 24 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=134870 $D=1
M136 260 24 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=139500 $D=1
M137 261 24 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=144130 $D=1
M138 9 25 262 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=134870 $D=1
M139 9 25 263 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=139500 $D=1
M140 9 25 264 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=144130 $D=1
M141 265 26 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=134870 $D=1
M142 266 26 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=139500 $D=1
M143 267 26 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=144130 $D=1
M144 268 25 223 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=134870 $D=1
M145 269 25 224 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=139500 $D=1
M146 270 25 225 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=144130 $D=1
M147 9 268 945 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=134870 $D=1
M148 9 269 946 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=139500 $D=1
M149 9 270 947 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=144130 $D=1
M150 271 945 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=134870 $D=1
M151 272 946 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=139500 $D=1
M152 273 947 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=144130 $D=1
M153 268 262 271 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=134870 $D=1
M154 269 263 272 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=139500 $D=1
M155 270 264 273 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=144130 $D=1
M156 271 26 238 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=134870 $D=1
M157 272 26 239 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=139500 $D=1
M158 273 26 240 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=144130 $D=1
M159 244 27 271 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=134870 $D=1
M160 245 27 272 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=139500 $D=1
M161 246 27 273 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=144130 $D=1
M162 274 27 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=134870 $D=1
M163 275 27 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=139500 $D=1
M164 276 27 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=144130 $D=1
M165 9 28 277 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=134870 $D=1
M166 9 28 278 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=139500 $D=1
M167 9 28 279 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=144130 $D=1
M168 280 29 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=134870 $D=1
M169 281 29 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=139500 $D=1
M170 282 29 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=144130 $D=1
M171 283 28 223 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=134870 $D=1
M172 284 28 224 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=139500 $D=1
M173 285 28 225 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=144130 $D=1
M174 9 283 948 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=134870 $D=1
M175 9 284 949 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=139500 $D=1
M176 9 285 950 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=144130 $D=1
M177 286 948 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=134870 $D=1
M178 287 949 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=139500 $D=1
M179 288 950 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=144130 $D=1
M180 283 277 286 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=134870 $D=1
M181 284 278 287 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=139500 $D=1
M182 285 279 288 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=144130 $D=1
M183 286 29 238 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=134870 $D=1
M184 287 29 239 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=139500 $D=1
M185 288 29 240 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=144130 $D=1
M186 244 30 286 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=134870 $D=1
M187 245 30 287 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=139500 $D=1
M188 246 30 288 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=144130 $D=1
M189 289 30 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=134870 $D=1
M190 290 30 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=139500 $D=1
M191 291 30 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=144130 $D=1
M192 9 31 292 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=134870 $D=1
M193 9 31 293 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=139500 $D=1
M194 9 31 294 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=144130 $D=1
M195 295 32 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=134870 $D=1
M196 296 32 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=139500 $D=1
M197 297 32 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=144130 $D=1
M198 298 31 223 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=134870 $D=1
M199 299 31 224 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=139500 $D=1
M200 300 31 225 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=144130 $D=1
M201 9 298 951 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=134870 $D=1
M202 9 299 952 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=139500 $D=1
M203 9 300 953 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=144130 $D=1
M204 301 951 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=134870 $D=1
M205 302 952 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=139500 $D=1
M206 303 953 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=144130 $D=1
M207 298 292 301 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=134870 $D=1
M208 299 293 302 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=139500 $D=1
M209 300 294 303 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=144130 $D=1
M210 301 32 238 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=134870 $D=1
M211 302 32 239 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=139500 $D=1
M212 303 32 240 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=144130 $D=1
M213 244 33 301 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=134870 $D=1
M214 245 33 302 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=139500 $D=1
M215 246 33 303 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=144130 $D=1
M216 304 33 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=134870 $D=1
M217 305 33 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=139500 $D=1
M218 306 33 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=144130 $D=1
M219 9 34 307 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=134870 $D=1
M220 9 34 308 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=139500 $D=1
M221 9 34 309 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=144130 $D=1
M222 310 35 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=134870 $D=1
M223 311 35 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=139500 $D=1
M224 312 35 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=144130 $D=1
M225 313 34 223 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=134870 $D=1
M226 314 34 224 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=139500 $D=1
M227 315 34 225 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=144130 $D=1
M228 9 313 954 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=134870 $D=1
M229 9 314 955 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=139500 $D=1
M230 9 315 956 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=144130 $D=1
M231 316 954 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=134870 $D=1
M232 317 955 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=139500 $D=1
M233 318 956 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=144130 $D=1
M234 313 307 316 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=134870 $D=1
M235 314 308 317 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=139500 $D=1
M236 315 309 318 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=144130 $D=1
M237 316 35 238 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=134870 $D=1
M238 317 35 239 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=139500 $D=1
M239 318 35 240 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=144130 $D=1
M240 244 36 316 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=134870 $D=1
M241 245 36 317 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=139500 $D=1
M242 246 36 318 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=144130 $D=1
M243 319 36 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=134870 $D=1
M244 320 36 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=139500 $D=1
M245 321 36 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=144130 $D=1
M246 9 37 322 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=134870 $D=1
M247 9 37 323 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=139500 $D=1
M248 9 37 324 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=144130 $D=1
M249 325 38 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=134870 $D=1
M250 326 38 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=139500 $D=1
M251 327 38 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=144130 $D=1
M252 328 37 223 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=134870 $D=1
M253 329 37 224 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=139500 $D=1
M254 330 37 225 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=144130 $D=1
M255 9 328 957 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=134870 $D=1
M256 9 329 958 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=139500 $D=1
M257 9 330 959 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=144130 $D=1
M258 331 957 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=134870 $D=1
M259 332 958 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=139500 $D=1
M260 333 959 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=144130 $D=1
M261 328 322 331 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=134870 $D=1
M262 329 323 332 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=139500 $D=1
M263 330 324 333 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=144130 $D=1
M264 331 38 238 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=134870 $D=1
M265 332 38 239 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=139500 $D=1
M266 333 38 240 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=144130 $D=1
M267 244 39 331 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=134870 $D=1
M268 245 39 332 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=139500 $D=1
M269 246 39 333 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=144130 $D=1
M270 334 39 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=134870 $D=1
M271 335 39 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=139500 $D=1
M272 336 39 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=144130 $D=1
M273 9 40 337 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=134870 $D=1
M274 9 40 338 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=139500 $D=1
M275 9 40 339 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=144130 $D=1
M276 340 41 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=134870 $D=1
M277 341 41 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=139500 $D=1
M278 342 41 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=144130 $D=1
M279 343 40 223 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=134870 $D=1
M280 344 40 224 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=139500 $D=1
M281 345 40 225 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=144130 $D=1
M282 9 343 960 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=134870 $D=1
M283 9 344 961 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=139500 $D=1
M284 9 345 962 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=144130 $D=1
M285 346 960 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=134870 $D=1
M286 347 961 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=139500 $D=1
M287 348 962 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=144130 $D=1
M288 343 337 346 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=134870 $D=1
M289 344 338 347 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=139500 $D=1
M290 345 339 348 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=144130 $D=1
M291 346 41 238 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=134870 $D=1
M292 347 41 239 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=139500 $D=1
M293 348 41 240 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=144130 $D=1
M294 244 42 346 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=134870 $D=1
M295 245 42 347 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=139500 $D=1
M296 246 42 348 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=144130 $D=1
M297 349 42 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=134870 $D=1
M298 350 42 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=139500 $D=1
M299 351 42 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=144130 $D=1
M300 9 43 352 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=134870 $D=1
M301 9 43 353 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=139500 $D=1
M302 9 43 354 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=144130 $D=1
M303 355 44 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=134870 $D=1
M304 356 44 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=139500 $D=1
M305 357 44 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=144130 $D=1
M306 358 43 223 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=134870 $D=1
M307 359 43 224 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=139500 $D=1
M308 360 43 225 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=144130 $D=1
M309 9 358 963 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=134870 $D=1
M310 9 359 964 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=139500 $D=1
M311 9 360 965 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=144130 $D=1
M312 361 963 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=134870 $D=1
M313 362 964 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=139500 $D=1
M314 363 965 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=144130 $D=1
M315 358 352 361 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=134870 $D=1
M316 359 353 362 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=139500 $D=1
M317 360 354 363 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=144130 $D=1
M318 361 44 238 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=134870 $D=1
M319 362 44 239 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=139500 $D=1
M320 363 44 240 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=144130 $D=1
M321 244 45 361 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=134870 $D=1
M322 245 45 362 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=139500 $D=1
M323 246 45 363 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=144130 $D=1
M324 364 45 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=134870 $D=1
M325 365 45 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=139500 $D=1
M326 366 45 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=144130 $D=1
M327 9 46 367 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=134870 $D=1
M328 9 46 368 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=139500 $D=1
M329 9 46 369 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=144130 $D=1
M330 370 47 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=134870 $D=1
M331 371 47 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=139500 $D=1
M332 372 47 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=144130 $D=1
M333 373 46 223 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=134870 $D=1
M334 374 46 224 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=139500 $D=1
M335 375 46 225 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=144130 $D=1
M336 9 373 966 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=134870 $D=1
M337 9 374 967 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=139500 $D=1
M338 9 375 968 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=144130 $D=1
M339 376 966 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=134870 $D=1
M340 377 967 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=139500 $D=1
M341 378 968 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=144130 $D=1
M342 373 367 376 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=134870 $D=1
M343 374 368 377 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=139500 $D=1
M344 375 369 378 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=144130 $D=1
M345 376 47 238 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=134870 $D=1
M346 377 47 239 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=139500 $D=1
M347 378 47 240 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=144130 $D=1
M348 244 48 376 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=134870 $D=1
M349 245 48 377 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=139500 $D=1
M350 246 48 378 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=144130 $D=1
M351 379 48 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=134870 $D=1
M352 380 48 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=139500 $D=1
M353 381 48 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=144130 $D=1
M354 9 49 382 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=134870 $D=1
M355 9 49 383 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=139500 $D=1
M356 9 49 384 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=144130 $D=1
M357 385 50 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=134870 $D=1
M358 386 50 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=139500 $D=1
M359 387 50 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=144130 $D=1
M360 388 49 223 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=134870 $D=1
M361 389 49 224 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=139500 $D=1
M362 390 49 225 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=144130 $D=1
M363 9 388 969 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=134870 $D=1
M364 9 389 970 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=139500 $D=1
M365 9 390 971 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=144130 $D=1
M366 391 969 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=134870 $D=1
M367 392 970 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=139500 $D=1
M368 393 971 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=144130 $D=1
M369 388 382 391 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=134870 $D=1
M370 389 383 392 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=139500 $D=1
M371 390 384 393 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=144130 $D=1
M372 391 50 238 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=134870 $D=1
M373 392 50 239 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=139500 $D=1
M374 393 50 240 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=144130 $D=1
M375 244 51 391 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=134870 $D=1
M376 245 51 392 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=139500 $D=1
M377 246 51 393 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=144130 $D=1
M378 394 51 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=134870 $D=1
M379 395 51 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=139500 $D=1
M380 396 51 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=144130 $D=1
M381 9 52 397 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=134870 $D=1
M382 9 52 398 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=139500 $D=1
M383 9 52 399 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=144130 $D=1
M384 400 53 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=134870 $D=1
M385 401 53 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=139500 $D=1
M386 402 53 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=144130 $D=1
M387 403 52 223 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=134870 $D=1
M388 404 52 224 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=139500 $D=1
M389 405 52 225 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=144130 $D=1
M390 9 403 972 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=134870 $D=1
M391 9 404 973 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=139500 $D=1
M392 9 405 974 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=144130 $D=1
M393 406 972 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=134870 $D=1
M394 407 973 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=139500 $D=1
M395 408 974 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=144130 $D=1
M396 403 397 406 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=134870 $D=1
M397 404 398 407 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=139500 $D=1
M398 405 399 408 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=144130 $D=1
M399 406 53 238 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=134870 $D=1
M400 407 53 239 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=139500 $D=1
M401 408 53 240 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=144130 $D=1
M402 244 54 406 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=134870 $D=1
M403 245 54 407 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=139500 $D=1
M404 246 54 408 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=144130 $D=1
M405 409 54 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=134870 $D=1
M406 410 54 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=139500 $D=1
M407 411 54 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=144130 $D=1
M408 9 55 412 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=134870 $D=1
M409 9 55 413 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=139500 $D=1
M410 9 55 414 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=144130 $D=1
M411 415 56 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=134870 $D=1
M412 416 56 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=139500 $D=1
M413 417 56 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=144130 $D=1
M414 418 55 223 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=134870 $D=1
M415 419 55 224 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=139500 $D=1
M416 420 55 225 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=144130 $D=1
M417 9 418 975 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=134870 $D=1
M418 9 419 976 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=139500 $D=1
M419 9 420 977 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=144130 $D=1
M420 421 975 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=134870 $D=1
M421 422 976 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=139500 $D=1
M422 423 977 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=144130 $D=1
M423 418 412 421 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=134870 $D=1
M424 419 413 422 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=139500 $D=1
M425 420 414 423 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=144130 $D=1
M426 421 56 238 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=134870 $D=1
M427 422 56 239 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=139500 $D=1
M428 423 56 240 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=144130 $D=1
M429 244 57 421 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=134870 $D=1
M430 245 57 422 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=139500 $D=1
M431 246 57 423 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=144130 $D=1
M432 424 57 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=134870 $D=1
M433 425 57 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=139500 $D=1
M434 426 57 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=144130 $D=1
M435 9 58 427 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=134870 $D=1
M436 9 58 428 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=139500 $D=1
M437 9 58 429 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=144130 $D=1
M438 430 59 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=134870 $D=1
M439 431 59 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=139500 $D=1
M440 432 59 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=144130 $D=1
M441 433 58 223 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=134870 $D=1
M442 434 58 224 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=139500 $D=1
M443 435 58 225 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=144130 $D=1
M444 9 433 978 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=134870 $D=1
M445 9 434 979 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=139500 $D=1
M446 9 435 980 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=144130 $D=1
M447 436 978 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=134870 $D=1
M448 437 979 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=139500 $D=1
M449 438 980 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=144130 $D=1
M450 433 427 436 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=134870 $D=1
M451 434 428 437 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=139500 $D=1
M452 435 429 438 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=144130 $D=1
M453 436 59 238 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=134870 $D=1
M454 437 59 239 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=139500 $D=1
M455 438 59 240 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=144130 $D=1
M456 244 60 436 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=134870 $D=1
M457 245 60 437 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=139500 $D=1
M458 246 60 438 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=144130 $D=1
M459 439 60 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=134870 $D=1
M460 440 60 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=139500 $D=1
M461 441 60 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=144130 $D=1
M462 9 61 442 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=134870 $D=1
M463 9 61 443 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=139500 $D=1
M464 9 61 444 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=144130 $D=1
M465 445 62 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=134870 $D=1
M466 446 62 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=139500 $D=1
M467 447 62 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=144130 $D=1
M468 448 61 223 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=134870 $D=1
M469 449 61 224 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=139500 $D=1
M470 450 61 225 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=144130 $D=1
M471 9 448 981 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=134870 $D=1
M472 9 449 982 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=139500 $D=1
M473 9 450 983 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=144130 $D=1
M474 451 981 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=134870 $D=1
M475 452 982 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=139500 $D=1
M476 453 983 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=144130 $D=1
M477 448 442 451 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=134870 $D=1
M478 449 443 452 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=139500 $D=1
M479 450 444 453 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=144130 $D=1
M480 451 62 238 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=134870 $D=1
M481 452 62 239 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=139500 $D=1
M482 453 62 240 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=144130 $D=1
M483 244 63 451 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=134870 $D=1
M484 245 63 452 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=139500 $D=1
M485 246 63 453 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=144130 $D=1
M486 454 63 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=134870 $D=1
M487 455 63 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=139500 $D=1
M488 456 63 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=144130 $D=1
M489 9 64 457 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=134870 $D=1
M490 9 64 458 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=139500 $D=1
M491 9 64 459 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=144130 $D=1
M492 460 65 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=134870 $D=1
M493 461 65 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=139500 $D=1
M494 462 65 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=144130 $D=1
M495 463 64 223 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=134870 $D=1
M496 464 64 224 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=139500 $D=1
M497 465 64 225 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=144130 $D=1
M498 9 463 984 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=134870 $D=1
M499 9 464 985 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=139500 $D=1
M500 9 465 986 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=144130 $D=1
M501 466 984 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=134870 $D=1
M502 467 985 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=139500 $D=1
M503 468 986 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=144130 $D=1
M504 463 457 466 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=134870 $D=1
M505 464 458 467 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=139500 $D=1
M506 465 459 468 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=144130 $D=1
M507 466 65 238 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=134870 $D=1
M508 467 65 239 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=139500 $D=1
M509 468 65 240 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=144130 $D=1
M510 244 66 466 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=134870 $D=1
M511 245 66 467 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=139500 $D=1
M512 246 66 468 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=144130 $D=1
M513 469 66 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=134870 $D=1
M514 470 66 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=139500 $D=1
M515 471 66 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=144130 $D=1
M516 9 67 472 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=134870 $D=1
M517 9 67 473 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=139500 $D=1
M518 9 67 474 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=144130 $D=1
M519 475 68 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=134870 $D=1
M520 476 68 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=139500 $D=1
M521 477 68 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=144130 $D=1
M522 478 67 223 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=134870 $D=1
M523 479 67 224 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=139500 $D=1
M524 480 67 225 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=144130 $D=1
M525 9 478 987 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=134870 $D=1
M526 9 479 988 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=139500 $D=1
M527 9 480 989 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=144130 $D=1
M528 481 987 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=134870 $D=1
M529 482 988 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=139500 $D=1
M530 483 989 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=144130 $D=1
M531 478 472 481 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=134870 $D=1
M532 479 473 482 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=139500 $D=1
M533 480 474 483 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=144130 $D=1
M534 481 68 238 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=134870 $D=1
M535 482 68 239 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=139500 $D=1
M536 483 68 240 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=144130 $D=1
M537 244 69 481 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=134870 $D=1
M538 245 69 482 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=139500 $D=1
M539 246 69 483 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=144130 $D=1
M540 484 69 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=134870 $D=1
M541 485 69 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=139500 $D=1
M542 486 69 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=144130 $D=1
M543 9 70 487 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=134870 $D=1
M544 9 70 488 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=139500 $D=1
M545 9 70 489 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=144130 $D=1
M546 490 71 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=134870 $D=1
M547 491 71 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=139500 $D=1
M548 492 71 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=144130 $D=1
M549 493 70 223 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=134870 $D=1
M550 494 70 224 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=139500 $D=1
M551 495 70 225 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=144130 $D=1
M552 9 493 990 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=134870 $D=1
M553 9 494 991 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=139500 $D=1
M554 9 495 992 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=144130 $D=1
M555 496 990 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=134870 $D=1
M556 497 991 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=139500 $D=1
M557 498 992 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=144130 $D=1
M558 493 487 496 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=134870 $D=1
M559 494 488 497 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=139500 $D=1
M560 495 489 498 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=144130 $D=1
M561 496 71 238 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=134870 $D=1
M562 497 71 239 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=139500 $D=1
M563 498 71 240 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=144130 $D=1
M564 244 72 496 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=134870 $D=1
M565 245 72 497 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=139500 $D=1
M566 246 72 498 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=144130 $D=1
M567 499 72 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=134870 $D=1
M568 500 72 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=139500 $D=1
M569 501 72 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=144130 $D=1
M570 9 73 502 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=134870 $D=1
M571 9 73 503 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=139500 $D=1
M572 9 73 504 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=144130 $D=1
M573 505 74 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=134870 $D=1
M574 506 74 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=139500 $D=1
M575 507 74 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=144130 $D=1
M576 508 73 223 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=134870 $D=1
M577 509 73 224 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=139500 $D=1
M578 510 73 225 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=144130 $D=1
M579 9 508 993 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=134870 $D=1
M580 9 509 994 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=139500 $D=1
M581 9 510 995 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=144130 $D=1
M582 511 993 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=134870 $D=1
M583 512 994 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=139500 $D=1
M584 513 995 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=144130 $D=1
M585 508 502 511 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=134870 $D=1
M586 509 503 512 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=139500 $D=1
M587 510 504 513 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=144130 $D=1
M588 511 74 238 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=134870 $D=1
M589 512 74 239 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=139500 $D=1
M590 513 74 240 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=144130 $D=1
M591 244 75 511 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=134870 $D=1
M592 245 75 512 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=139500 $D=1
M593 246 75 513 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=144130 $D=1
M594 514 75 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=134870 $D=1
M595 515 75 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=139500 $D=1
M596 516 75 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=144130 $D=1
M597 9 76 517 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=134870 $D=1
M598 9 76 518 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=139500 $D=1
M599 9 76 519 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=144130 $D=1
M600 520 77 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=134870 $D=1
M601 521 77 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=139500 $D=1
M602 522 77 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=144130 $D=1
M603 523 76 223 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=134870 $D=1
M604 524 76 224 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=139500 $D=1
M605 525 76 225 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=144130 $D=1
M606 9 523 996 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=134870 $D=1
M607 9 524 997 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=139500 $D=1
M608 9 525 998 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=144130 $D=1
M609 526 996 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=134870 $D=1
M610 527 997 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=139500 $D=1
M611 528 998 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=144130 $D=1
M612 523 517 526 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=134870 $D=1
M613 524 518 527 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=139500 $D=1
M614 525 519 528 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=144130 $D=1
M615 526 77 238 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=134870 $D=1
M616 527 77 239 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=139500 $D=1
M617 528 77 240 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=144130 $D=1
M618 244 78 526 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=134870 $D=1
M619 245 78 527 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=139500 $D=1
M620 246 78 528 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=144130 $D=1
M621 529 78 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=134870 $D=1
M622 530 78 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=139500 $D=1
M623 531 78 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=144130 $D=1
M624 9 79 532 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=134870 $D=1
M625 9 79 533 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=139500 $D=1
M626 9 79 534 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=144130 $D=1
M627 535 80 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=134870 $D=1
M628 536 80 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=139500 $D=1
M629 537 80 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=144130 $D=1
M630 538 79 223 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=134870 $D=1
M631 539 79 224 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=139500 $D=1
M632 540 79 225 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=144130 $D=1
M633 9 538 999 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=134870 $D=1
M634 9 539 1000 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=139500 $D=1
M635 9 540 1001 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=144130 $D=1
M636 541 999 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=134870 $D=1
M637 542 1000 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=139500 $D=1
M638 543 1001 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=144130 $D=1
M639 538 532 541 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=134870 $D=1
M640 539 533 542 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=139500 $D=1
M641 540 534 543 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=144130 $D=1
M642 541 80 238 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=134870 $D=1
M643 542 80 239 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=139500 $D=1
M644 543 80 240 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=144130 $D=1
M645 244 81 541 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=134870 $D=1
M646 245 81 542 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=139500 $D=1
M647 246 81 543 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=144130 $D=1
M648 544 81 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=134870 $D=1
M649 545 81 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=139500 $D=1
M650 546 81 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=144130 $D=1
M651 9 82 547 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=134870 $D=1
M652 9 82 548 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=139500 $D=1
M653 9 82 549 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=144130 $D=1
M654 550 83 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=134870 $D=1
M655 551 83 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=139500 $D=1
M656 552 83 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=144130 $D=1
M657 553 82 223 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=134870 $D=1
M658 554 82 224 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=139500 $D=1
M659 555 82 225 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=144130 $D=1
M660 9 553 1002 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=134870 $D=1
M661 9 554 1003 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=139500 $D=1
M662 9 555 1004 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=144130 $D=1
M663 556 1002 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=134870 $D=1
M664 557 1003 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=139500 $D=1
M665 558 1004 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=144130 $D=1
M666 553 547 556 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=134870 $D=1
M667 554 548 557 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=139500 $D=1
M668 555 549 558 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=144130 $D=1
M669 556 83 238 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=134870 $D=1
M670 557 83 239 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=139500 $D=1
M671 558 83 240 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=144130 $D=1
M672 244 84 556 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=134870 $D=1
M673 245 84 557 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=139500 $D=1
M674 246 84 558 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=144130 $D=1
M675 559 84 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=134870 $D=1
M676 560 84 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=139500 $D=1
M677 561 84 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=144130 $D=1
M678 9 85 562 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=134870 $D=1
M679 9 85 563 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=139500 $D=1
M680 9 85 564 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=144130 $D=1
M681 565 86 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=134870 $D=1
M682 566 86 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=139500 $D=1
M683 567 86 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=144130 $D=1
M684 568 85 223 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=134870 $D=1
M685 569 85 224 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=139500 $D=1
M686 570 85 225 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=144130 $D=1
M687 9 568 1005 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=134870 $D=1
M688 9 569 1006 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=139500 $D=1
M689 9 570 1007 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=144130 $D=1
M690 571 1005 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=134870 $D=1
M691 572 1006 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=139500 $D=1
M692 573 1007 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=144130 $D=1
M693 568 562 571 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=134870 $D=1
M694 569 563 572 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=139500 $D=1
M695 570 564 573 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=144130 $D=1
M696 571 86 238 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=134870 $D=1
M697 572 86 239 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=139500 $D=1
M698 573 86 240 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=144130 $D=1
M699 244 87 571 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=134870 $D=1
M700 245 87 572 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=139500 $D=1
M701 246 87 573 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=144130 $D=1
M702 574 87 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=134870 $D=1
M703 575 87 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=139500 $D=1
M704 576 87 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=144130 $D=1
M705 9 88 577 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=134870 $D=1
M706 9 88 578 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=139500 $D=1
M707 9 88 579 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=144130 $D=1
M708 580 89 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=134870 $D=1
M709 581 89 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=139500 $D=1
M710 582 89 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=144130 $D=1
M711 583 88 223 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=134870 $D=1
M712 584 88 224 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=139500 $D=1
M713 585 88 225 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=144130 $D=1
M714 9 583 1008 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=134870 $D=1
M715 9 584 1009 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=139500 $D=1
M716 9 585 1010 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=144130 $D=1
M717 586 1008 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=134870 $D=1
M718 587 1009 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=139500 $D=1
M719 588 1010 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=144130 $D=1
M720 583 577 586 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=134870 $D=1
M721 584 578 587 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=139500 $D=1
M722 585 579 588 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=144130 $D=1
M723 586 89 238 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=134870 $D=1
M724 587 89 239 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=139500 $D=1
M725 588 89 240 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=144130 $D=1
M726 244 90 586 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=134870 $D=1
M727 245 90 587 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=139500 $D=1
M728 246 90 588 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=144130 $D=1
M729 589 90 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=134870 $D=1
M730 590 90 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=139500 $D=1
M731 591 90 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=144130 $D=1
M732 9 91 592 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=134870 $D=1
M733 9 91 593 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=139500 $D=1
M734 9 91 594 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=144130 $D=1
M735 595 92 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=134870 $D=1
M736 596 92 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=139500 $D=1
M737 597 92 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=144130 $D=1
M738 598 91 223 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=134870 $D=1
M739 599 91 224 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=139500 $D=1
M740 600 91 225 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=144130 $D=1
M741 9 598 1011 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=134870 $D=1
M742 9 599 1012 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=139500 $D=1
M743 9 600 1013 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=144130 $D=1
M744 601 1011 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=134870 $D=1
M745 602 1012 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=139500 $D=1
M746 603 1013 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=144130 $D=1
M747 598 592 601 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=134870 $D=1
M748 599 593 602 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=139500 $D=1
M749 600 594 603 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=144130 $D=1
M750 601 92 238 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=134870 $D=1
M751 602 92 239 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=139500 $D=1
M752 603 92 240 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=144130 $D=1
M753 244 93 601 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=134870 $D=1
M754 245 93 602 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=139500 $D=1
M755 246 93 603 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=144130 $D=1
M756 604 93 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=134870 $D=1
M757 605 93 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=139500 $D=1
M758 606 93 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=144130 $D=1
M759 9 94 607 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=134870 $D=1
M760 9 94 608 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=139500 $D=1
M761 9 94 609 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=144130 $D=1
M762 610 95 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=134870 $D=1
M763 611 95 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=139500 $D=1
M764 612 95 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=144130 $D=1
M765 613 94 223 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=134870 $D=1
M766 614 94 224 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=139500 $D=1
M767 615 94 225 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=144130 $D=1
M768 9 613 1014 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=134870 $D=1
M769 9 614 1015 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=139500 $D=1
M770 9 615 1016 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=144130 $D=1
M771 616 1014 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=134870 $D=1
M772 617 1015 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=139500 $D=1
M773 618 1016 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=144130 $D=1
M774 613 607 616 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=134870 $D=1
M775 614 608 617 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=139500 $D=1
M776 615 609 618 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=144130 $D=1
M777 616 95 238 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=134870 $D=1
M778 617 95 239 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=139500 $D=1
M779 618 95 240 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=144130 $D=1
M780 244 96 616 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=134870 $D=1
M781 245 96 617 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=139500 $D=1
M782 246 96 618 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=144130 $D=1
M783 619 96 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=134870 $D=1
M784 620 96 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=139500 $D=1
M785 621 96 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=144130 $D=1
M786 9 97 622 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=134870 $D=1
M787 9 97 623 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=139500 $D=1
M788 9 97 624 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=144130 $D=1
M789 625 98 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=134870 $D=1
M790 626 98 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=139500 $D=1
M791 627 98 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=144130 $D=1
M792 628 97 223 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=134870 $D=1
M793 629 97 224 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=139500 $D=1
M794 630 97 225 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=144130 $D=1
M795 9 628 1017 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=134870 $D=1
M796 9 629 1018 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=139500 $D=1
M797 9 630 1019 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=144130 $D=1
M798 631 1017 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=134870 $D=1
M799 632 1018 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=139500 $D=1
M800 633 1019 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=144130 $D=1
M801 628 622 631 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=134870 $D=1
M802 629 623 632 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=139500 $D=1
M803 630 624 633 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=144130 $D=1
M804 631 98 238 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=134870 $D=1
M805 632 98 239 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=139500 $D=1
M806 633 98 240 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=144130 $D=1
M807 244 99 631 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=134870 $D=1
M808 245 99 632 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=139500 $D=1
M809 246 99 633 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=144130 $D=1
M810 634 99 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=134870 $D=1
M811 635 99 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=139500 $D=1
M812 636 99 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=144130 $D=1
M813 9 100 637 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=134870 $D=1
M814 9 100 638 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=139500 $D=1
M815 9 100 639 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=144130 $D=1
M816 640 101 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=134870 $D=1
M817 641 101 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=139500 $D=1
M818 642 101 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=144130 $D=1
M819 643 100 223 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=134870 $D=1
M820 644 100 224 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=139500 $D=1
M821 645 100 225 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=144130 $D=1
M822 9 643 1020 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=134870 $D=1
M823 9 644 1021 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=139500 $D=1
M824 9 645 1022 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=144130 $D=1
M825 646 1020 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=134870 $D=1
M826 647 1021 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=139500 $D=1
M827 648 1022 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=144130 $D=1
M828 643 637 646 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=134870 $D=1
M829 644 638 647 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=139500 $D=1
M830 645 639 648 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=144130 $D=1
M831 646 101 238 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=134870 $D=1
M832 647 101 239 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=139500 $D=1
M833 648 101 240 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=144130 $D=1
M834 244 102 646 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=134870 $D=1
M835 245 102 647 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=139500 $D=1
M836 246 102 648 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=144130 $D=1
M837 649 102 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=134870 $D=1
M838 650 102 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=139500 $D=1
M839 651 102 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=144130 $D=1
M840 9 103 652 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=134870 $D=1
M841 9 103 653 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=139500 $D=1
M842 9 103 654 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=144130 $D=1
M843 655 104 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=134870 $D=1
M844 656 104 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=139500 $D=1
M845 657 104 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=144130 $D=1
M846 658 103 223 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=134870 $D=1
M847 659 103 224 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=139500 $D=1
M848 660 103 225 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=144130 $D=1
M849 9 658 1023 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=134870 $D=1
M850 9 659 1024 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=139500 $D=1
M851 9 660 1025 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=144130 $D=1
M852 661 1023 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=134870 $D=1
M853 662 1024 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=139500 $D=1
M854 663 1025 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=144130 $D=1
M855 658 652 661 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=134870 $D=1
M856 659 653 662 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=139500 $D=1
M857 660 654 663 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=144130 $D=1
M858 661 104 238 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=134870 $D=1
M859 662 104 239 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=139500 $D=1
M860 663 104 240 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=144130 $D=1
M861 244 105 661 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=134870 $D=1
M862 245 105 662 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=139500 $D=1
M863 246 105 663 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=144130 $D=1
M864 664 105 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=134870 $D=1
M865 665 105 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=139500 $D=1
M866 666 105 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=144130 $D=1
M867 9 106 667 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=134870 $D=1
M868 9 106 668 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=139500 $D=1
M869 9 106 669 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=144130 $D=1
M870 670 107 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=134870 $D=1
M871 671 107 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=139500 $D=1
M872 672 107 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=144130 $D=1
M873 673 106 223 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=134870 $D=1
M874 674 106 224 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=139500 $D=1
M875 675 106 225 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=144130 $D=1
M876 9 673 1026 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=134870 $D=1
M877 9 674 1027 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=139500 $D=1
M878 9 675 1028 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=144130 $D=1
M879 676 1026 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=134870 $D=1
M880 677 1027 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=139500 $D=1
M881 678 1028 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=144130 $D=1
M882 673 667 676 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=134870 $D=1
M883 674 668 677 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=139500 $D=1
M884 675 669 678 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=144130 $D=1
M885 676 107 238 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=134870 $D=1
M886 677 107 239 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=139500 $D=1
M887 678 107 240 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=144130 $D=1
M888 244 108 676 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=134870 $D=1
M889 245 108 677 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=139500 $D=1
M890 246 108 678 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=144130 $D=1
M891 679 108 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=134870 $D=1
M892 680 108 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=139500 $D=1
M893 681 108 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=144130 $D=1
M894 9 109 682 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=134870 $D=1
M895 9 109 683 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=139500 $D=1
M896 9 109 684 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=144130 $D=1
M897 685 110 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=134870 $D=1
M898 686 110 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=139500 $D=1
M899 687 110 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=144130 $D=1
M900 688 109 223 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=134870 $D=1
M901 689 109 224 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=139500 $D=1
M902 690 109 225 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=144130 $D=1
M903 9 688 1029 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=134870 $D=1
M904 9 689 1030 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=139500 $D=1
M905 9 690 1031 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=144130 $D=1
M906 691 1029 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=134870 $D=1
M907 692 1030 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=139500 $D=1
M908 693 1031 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=144130 $D=1
M909 688 682 691 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=134870 $D=1
M910 689 683 692 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=139500 $D=1
M911 690 684 693 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=144130 $D=1
M912 691 110 238 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=134870 $D=1
M913 692 110 239 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=139500 $D=1
M914 693 110 240 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=144130 $D=1
M915 244 111 691 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=134870 $D=1
M916 245 111 692 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=139500 $D=1
M917 246 111 693 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=144130 $D=1
M918 694 111 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=134870 $D=1
M919 695 111 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=139500 $D=1
M920 696 111 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=144130 $D=1
M921 9 112 697 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=134870 $D=1
M922 9 112 698 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=139500 $D=1
M923 9 112 699 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=144130 $D=1
M924 700 113 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=134870 $D=1
M925 701 113 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=139500 $D=1
M926 702 113 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=144130 $D=1
M927 9 113 238 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=134870 $D=1
M928 9 113 239 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=139500 $D=1
M929 9 113 240 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=144130 $D=1
M930 244 112 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=134870 $D=1
M931 245 112 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=139500 $D=1
M932 246 112 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=144130 $D=1
M933 9 706 703 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=134870 $D=1
M934 9 707 704 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=139500 $D=1
M935 9 708 705 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=144130 $D=1
M936 706 114 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=134870 $D=1
M937 707 114 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=139500 $D=1
M938 708 114 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=144130 $D=1
M939 1032 238 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=134870 $D=1
M940 1033 239 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=139500 $D=1
M941 1034 240 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=144130 $D=1
M942 709 703 1032 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=134870 $D=1
M943 710 704 1033 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=139500 $D=1
M944 711 705 1034 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=144130 $D=1
M945 9 709 712 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=134870 $D=1
M946 9 710 713 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=139500 $D=1
M947 9 711 714 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=144130 $D=1
M948 1035 712 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=134870 $D=1
M949 1036 713 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=139500 $D=1
M950 1037 714 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=144130 $D=1
M951 709 706 1035 9 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=134870 $D=1
M952 710 707 1036 9 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=139500 $D=1
M953 711 708 1037 9 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=144130 $D=1
M954 9 718 715 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=134870 $D=1
M955 9 719 716 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=139500 $D=1
M956 9 720 717 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=144130 $D=1
M957 718 114 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=134870 $D=1
M958 719 114 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=139500 $D=1
M959 720 114 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=144130 $D=1
M960 1038 244 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=134870 $D=1
M961 1039 245 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=139500 $D=1
M962 1040 246 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=144130 $D=1
M963 721 715 1038 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=134870 $D=1
M964 722 716 1039 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=139500 $D=1
M965 723 717 1040 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=144130 $D=1
M966 9 721 115 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=134870 $D=1
M967 9 722 116 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=139500 $D=1
M968 9 723 117 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=144130 $D=1
M969 1041 115 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=134870 $D=1
M970 1042 116 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=139500 $D=1
M971 1043 117 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=144130 $D=1
M972 721 718 1041 9 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=134870 $D=1
M973 722 719 1042 9 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=139500 $D=1
M974 723 720 1043 9 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=144130 $D=1
M975 724 118 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=134870 $D=1
M976 725 118 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=139500 $D=1
M977 726 118 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=144130 $D=1
M978 727 724 712 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=134870 $D=1
M979 728 725 713 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=139500 $D=1
M980 729 726 714 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=144130 $D=1
M981 119 118 727 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=134870 $D=1
M982 120 118 728 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=139500 $D=1
M983 121 118 729 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=144130 $D=1
M984 730 122 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=134870 $D=1
M985 731 122 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=139500 $D=1
M986 732 122 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=144130 $D=1
M987 733 730 115 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=134870 $D=1
M988 734 731 116 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=139500 $D=1
M989 735 732 117 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=144130 $D=1
M990 1044 122 733 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=134870 $D=1
M991 1045 122 734 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=139500 $D=1
M992 1046 122 735 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=144130 $D=1
M993 9 115 1044 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=134870 $D=1
M994 9 116 1045 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=139500 $D=1
M995 9 117 1046 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=144130 $D=1
M996 736 123 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=134870 $D=1
M997 737 123 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=139500 $D=1
M998 738 123 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=144130 $D=1
M999 124 736 733 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=134870 $D=1
M1000 125 737 734 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=139500 $D=1
M1001 126 738 735 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=144130 $D=1
M1002 11 123 124 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=134870 $D=1
M1003 12 123 125 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=139500 $D=1
M1004 13 123 126 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=144130 $D=1
M1005 741 739 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=134870 $D=1
M1006 742 740 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=139500 $D=1
M1007 743 127 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=144130 $D=1
M1008 9 747 744 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=134870 $D=1
M1009 9 748 745 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=139500 $D=1
M1010 9 749 746 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=144130 $D=1
M1011 750 727 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=134870 $D=1
M1012 751 728 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=139500 $D=1
M1013 752 729 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=144130 $D=1
M1014 747 750 739 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=134870 $D=1
M1015 748 751 740 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=139500 $D=1
M1016 749 752 127 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=144130 $D=1
M1017 741 727 747 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=134870 $D=1
M1018 742 728 748 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=139500 $D=1
M1019 743 729 749 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=144130 $D=1
M1020 753 744 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=134870 $D=1
M1021 754 745 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=139500 $D=1
M1022 755 746 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=144130 $D=1
M1023 128 753 124 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=134870 $D=1
M1024 739 754 125 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=139500 $D=1
M1025 740 755 126 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=144130 $D=1
M1026 727 744 128 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=134870 $D=1
M1027 728 745 739 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=139500 $D=1
M1028 729 746 740 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=144130 $D=1
M1029 756 128 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=134870 $D=1
M1030 757 739 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=139500 $D=1
M1031 758 740 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=144130 $D=1
M1032 759 744 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=134870 $D=1
M1033 760 745 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=139500 $D=1
M1034 761 746 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=144130 $D=1
M1035 762 759 756 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=134870 $D=1
M1036 763 760 757 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=139500 $D=1
M1037 764 761 758 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=144130 $D=1
M1038 124 744 762 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=134870 $D=1
M1039 125 745 763 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=139500 $D=1
M1040 126 746 764 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=144130 $D=1
M1041 765 727 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=134870 $D=1
M1042 766 728 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=139500 $D=1
M1043 767 729 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=144130 $D=1
M1044 9 124 765 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=134870 $D=1
M1045 9 125 766 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=139500 $D=1
M1046 9 126 767 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=144130 $D=1
M1047 768 762 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=134870 $D=1
M1048 769 763 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=139500 $D=1
M1049 770 764 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=144130 $D=1
M1050 1074 727 9 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=134870 $D=1
M1051 1075 728 9 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=139500 $D=1
M1052 1076 729 9 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=144130 $D=1
M1053 771 124 1074 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=134870 $D=1
M1054 772 125 1075 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=139500 $D=1
M1055 773 126 1076 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=144130 $D=1
M1056 1077 727 9 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=134870 $D=1
M1057 1078 728 9 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=139500 $D=1
M1058 1079 729 9 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=144130 $D=1
M1059 774 124 1077 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=134870 $D=1
M1060 775 125 1078 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=139500 $D=1
M1061 776 126 1079 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=144130 $D=1
M1062 780 727 777 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=134870 $D=1
M1063 781 728 778 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=139500 $D=1
M1064 782 729 779 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=144130 $D=1
M1065 777 124 780 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=134870 $D=1
M1066 778 125 781 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=139500 $D=1
M1067 779 126 782 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=144130 $D=1
M1068 9 774 777 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=134870 $D=1
M1069 9 775 778 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=139500 $D=1
M1070 9 776 779 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=144130 $D=1
M1071 783 135 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=134870 $D=1
M1072 784 135 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=139500 $D=1
M1073 785 135 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=144130 $D=1
M1074 786 783 765 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=134870 $D=1
M1075 787 784 766 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=139500 $D=1
M1076 788 785 767 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=144130 $D=1
M1077 771 135 786 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=134870 $D=1
M1078 772 135 787 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=139500 $D=1
M1079 773 135 788 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=144130 $D=1
M1080 789 783 768 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=134870 $D=1
M1081 790 784 769 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=139500 $D=1
M1082 791 785 770 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=144130 $D=1
M1083 780 135 789 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=134870 $D=1
M1084 781 135 790 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=139500 $D=1
M1085 782 135 791 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=144130 $D=1
M1086 792 136 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=134870 $D=1
M1087 793 136 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=139500 $D=1
M1088 794 136 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=144130 $D=1
M1089 795 792 789 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=134870 $D=1
M1090 796 793 790 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=139500 $D=1
M1091 797 794 791 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=144130 $D=1
M1092 786 136 795 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=134870 $D=1
M1093 787 136 796 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=139500 $D=1
M1094 788 136 797 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=144130 $D=1
M1095 14 795 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=134870 $D=1
M1096 15 796 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=139500 $D=1
M1097 16 797 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=144130 $D=1
M1098 798 137 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=134870 $D=1
M1099 799 137 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=139500 $D=1
M1100 800 137 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=144130 $D=1
M1101 803 798 801 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=134870 $D=1
M1102 804 799 802 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=139500 $D=1
M1103 805 800 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=144130 $D=1
M1104 138 137 803 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=134870 $D=1
M1105 139 137 804 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=139500 $D=1
M1106 801 137 805 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=144130 $D=1
M1107 806 137 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=134870 $D=1
M1108 807 137 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=139500 $D=1
M1109 808 137 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=144130 $D=1
M1110 810 806 809 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=134870 $D=1
M1111 811 807 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=139500 $D=1
M1112 812 808 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=144130 $D=1
M1113 140 137 810 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=134870 $D=1
M1114 141 137 811 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=139500 $D=1
M1115 142 137 812 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=144130 $D=1
M1116 813 137 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=134870 $D=1
M1117 814 137 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=139500 $D=1
M1118 815 137 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=144130 $D=1
M1119 816 813 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=134870 $D=1
M1120 817 814 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=139500 $D=1
M1121 818 815 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=144130 $D=1
M1122 143 137 816 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=134870 $D=1
M1123 144 137 817 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=139500 $D=1
M1124 145 137 818 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=144130 $D=1
M1125 819 137 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=134870 $D=1
M1126 820 137 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=139500 $D=1
M1127 821 137 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=144130 $D=1
M1128 822 819 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=134870 $D=1
M1129 823 820 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=139500 $D=1
M1130 824 821 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=144130 $D=1
M1131 146 137 822 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=134870 $D=1
M1132 147 137 823 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=139500 $D=1
M1133 148 137 824 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=144130 $D=1
M1134 825 137 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=134870 $D=1
M1135 826 137 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=139500 $D=1
M1136 827 137 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=144130 $D=1
M1137 828 825 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=134870 $D=1
M1138 829 826 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=139500 $D=1
M1139 830 827 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=144130 $D=1
M1140 149 137 828 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=134870 $D=1
M1141 150 137 829 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=139500 $D=1
M1142 151 137 830 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=144130 $D=1
M1143 9 727 1047 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=134870 $D=1
M1144 9 728 1048 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=139500 $D=1
M1145 9 729 1049 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=144130 $D=1
M1146 139 1047 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=134870 $D=1
M1147 801 1048 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=139500 $D=1
M1148 802 1049 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=144130 $D=1
M1149 831 126 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=134870 $D=1
M1150 832 126 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=139500 $D=1
M1151 833 126 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=144130 $D=1
M1152 142 831 139 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=134870 $D=1
M1153 152 832 801 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=139500 $D=1
M1154 809 833 802 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=144130 $D=1
M1155 803 126 142 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=134870 $D=1
M1156 804 126 152 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=139500 $D=1
M1157 805 126 809 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=144130 $D=1
M1158 834 125 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=134870 $D=1
M1159 835 125 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=139500 $D=1
M1160 836 125 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=144130 $D=1
M1161 134 834 142 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=134870 $D=1
M1162 133 835 152 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=139500 $D=1
M1163 132 836 809 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=144130 $D=1
M1164 810 125 134 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=134870 $D=1
M1165 811 125 133 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=139500 $D=1
M1166 812 125 132 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=144130 $D=1
M1167 837 124 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=134870 $D=1
M1168 838 124 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=139500 $D=1
M1169 839 124 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=144130 $D=1
M1170 129 837 134 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=134870 $D=1
M1171 130 838 133 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=139500 $D=1
M1172 131 839 132 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=144130 $D=1
M1173 816 124 129 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=134870 $D=1
M1174 817 124 130 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=139500 $D=1
M1175 818 124 131 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=144130 $D=1
M1176 840 153 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=134870 $D=1
M1177 841 153 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=139500 $D=1
M1178 842 153 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=144130 $D=1
M1179 154 840 129 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=134870 $D=1
M1180 155 841 130 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=139500 $D=1
M1181 156 842 131 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=144130 $D=1
M1182 822 153 154 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=134870 $D=1
M1183 823 153 155 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=139500 $D=1
M1184 824 153 156 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=144130 $D=1
M1185 843 157 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=134870 $D=1
M1186 844 157 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=139500 $D=1
M1187 845 157 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=144130 $D=1
M1188 202 843 154 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=134870 $D=1
M1189 203 844 155 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=139500 $D=1
M1190 204 845 156 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=144130 $D=1
M1191 828 157 202 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=134870 $D=1
M1192 829 157 203 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=139500 $D=1
M1193 830 157 204 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=144130 $D=1
M1194 846 158 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=134870 $D=1
M1195 847 158 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=139500 $D=1
M1196 848 158 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=144130 $D=1
M1197 849 846 115 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=134870 $D=1
M1198 850 847 116 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=139500 $D=1
M1199 851 848 117 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=144130 $D=1
M1200 11 158 849 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=134870 $D=1
M1201 12 158 850 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=139500 $D=1
M1202 13 158 851 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=144130 $D=1
M1203 1080 712 9 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=134870 $D=1
M1204 1081 713 9 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=139500 $D=1
M1205 1082 714 9 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=144130 $D=1
M1206 852 849 1080 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=134870 $D=1
M1207 853 850 1081 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=139500 $D=1
M1208 854 851 1082 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=144130 $D=1
M1209 858 712 855 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=134870 $D=1
M1210 859 713 856 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=139500 $D=1
M1211 860 714 857 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=144130 $D=1
M1212 855 849 858 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=134870 $D=1
M1213 856 850 859 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=139500 $D=1
M1214 857 851 860 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=144130 $D=1
M1215 9 852 855 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=134870 $D=1
M1216 9 853 856 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=139500 $D=1
M1217 9 854 857 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=144130 $D=1
M1218 1083 159 9 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=134870 $D=1
M1219 1084 861 9 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=139500 $D=1
M1220 1085 862 9 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=144130 $D=1
M1221 1050 858 1083 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=134870 $D=1
M1222 1051 859 1084 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=139500 $D=1
M1223 1052 860 1085 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=144130 $D=1
M1224 861 1050 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=134870 $D=1
M1225 862 1051 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=139500 $D=1
M1226 160 1052 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=144130 $D=1
M1227 863 712 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=134870 $D=1
M1228 864 713 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=139500 $D=1
M1229 865 714 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=144130 $D=1
M1230 9 866 863 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=134870 $D=1
M1231 9 867 864 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=139500 $D=1
M1232 9 868 865 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=144130 $D=1
M1233 866 849 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=134870 $D=1
M1234 867 850 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=139500 $D=1
M1235 868 851 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=144130 $D=1
M1236 1086 863 9 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=134870 $D=1
M1237 1087 864 9 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=139500 $D=1
M1238 1088 865 9 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=144130 $D=1
M1239 869 159 1086 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=134870 $D=1
M1240 870 861 1087 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=139500 $D=1
M1241 871 862 1088 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=144130 $D=1
M1242 874 161 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=134870 $D=1
M1243 875 872 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=139500 $D=1
M1244 876 873 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=144130 $D=1
M1245 1089 869 9 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=134870 $D=1
M1246 1090 870 9 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=139500 $D=1
M1247 1091 871 9 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=144130 $D=1
M1248 872 874 1089 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=134870 $D=1
M1249 873 875 1090 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=139500 $D=1
M1250 162 876 1091 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=144130 $D=1
M1251 879 877 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=134870 $D=1
M1252 880 878 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=139500 $D=1
M1253 881 9 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=144130 $D=1
M1254 9 885 882 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=134870 $D=1
M1255 9 886 883 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=139500 $D=1
M1256 9 887 884 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=144130 $D=1
M1257 888 119 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=134870 $D=1
M1258 889 120 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=139500 $D=1
M1259 890 121 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=144130 $D=1
M1260 885 888 877 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=134870 $D=1
M1261 886 889 878 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=139500 $D=1
M1262 887 890 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=144130 $D=1
M1263 879 119 885 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=134870 $D=1
M1264 880 120 886 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=139500 $D=1
M1265 881 121 887 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=144130 $D=1
M1266 891 882 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=134870 $D=1
M1267 892 883 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=139500 $D=1
M1268 893 884 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=144130 $D=1
M1269 163 891 7 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=134870 $D=1
M1270 877 892 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=139500 $D=1
M1271 878 893 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=144130 $D=1
M1272 119 882 163 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=134870 $D=1
M1273 120 883 877 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=139500 $D=1
M1274 121 884 878 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=144130 $D=1
M1275 894 163 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=134870 $D=1
M1276 895 877 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=139500 $D=1
M1277 896 878 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=144130 $D=1
M1278 897 882 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=134870 $D=1
M1279 898 883 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=139500 $D=1
M1280 899 884 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=144130 $D=1
M1281 205 897 894 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=134870 $D=1
M1282 206 898 895 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=139500 $D=1
M1283 207 899 896 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=144130 $D=1
M1284 7 882 205 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=134870 $D=1
M1285 9 883 206 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=139500 $D=1
M1286 9 884 207 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=144130 $D=1
M1287 900 164 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=134870 $D=1
M1288 901 164 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=139500 $D=1
M1289 902 164 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=144130 $D=1
M1290 903 900 205 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=134870 $D=1
M1291 904 901 206 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=139500 $D=1
M1292 905 902 207 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=144130 $D=1
M1293 14 164 903 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=134870 $D=1
M1294 15 164 904 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=139500 $D=1
M1295 16 164 905 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=144130 $D=1
M1296 906 165 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=134870 $D=1
M1297 907 165 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=139500 $D=1
M1298 908 165 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=144130 $D=1
M1299 909 906 903 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=134870 $D=1
M1300 910 907 904 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=139500 $D=1
M1301 911 908 905 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=144130 $D=1
M1302 9 165 909 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=134870 $D=1
M1303 9 165 910 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=139500 $D=1
M1304 9 165 911 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=144130 $D=1
M1305 912 114 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=134870 $D=1
M1306 913 114 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=139500 $D=1
M1307 914 114 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=144130 $D=1
M1308 9 912 915 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=134870 $D=1
M1309 9 913 916 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=139500 $D=1
M1310 9 914 917 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=144130 $D=1
M1311 918 114 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=134870 $D=1
M1312 919 114 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=139500 $D=1
M1313 920 114 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=144130 $D=1
M1314 921 912 909 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=134870 $D=1
M1315 922 913 910 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=139500 $D=1
M1316 923 914 911 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=144130 $D=1
M1317 9 921 1053 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=134870 $D=1
M1318 9 922 1054 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=139500 $D=1
M1319 9 923 1055 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=144130 $D=1
M1320 924 1053 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=134870 $D=1
M1321 925 1054 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=139500 $D=1
M1322 926 1055 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=144130 $D=1
M1323 921 915 924 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=134870 $D=1
M1324 922 916 925 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=139500 $D=1
M1325 923 917 926 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=144130 $D=1
M1326 927 114 924 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=134870 $D=1
M1327 928 114 925 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=139500 $D=1
M1328 929 114 926 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=144130 $D=1
M1329 9 933 930 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=134870 $D=1
M1330 9 934 931 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=139500 $D=1
M1331 9 935 932 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=144130 $D=1
M1332 933 114 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=134870 $D=1
M1333 934 114 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=139500 $D=1
M1334 935 114 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=144130 $D=1
M1335 1056 927 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=134870 $D=1
M1336 1057 928 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=139500 $D=1
M1337 1058 929 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=144130 $D=1
M1338 936 930 1056 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=134870 $D=1
M1339 937 931 1057 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=139500 $D=1
M1340 938 932 1058 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=144130 $D=1
M1341 9 936 119 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=134870 $D=1
M1342 9 937 120 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=139500 $D=1
M1343 9 938 121 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=144130 $D=1
M1344 1059 119 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=134870 $D=1
M1345 1060 120 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=139500 $D=1
M1346 1061 121 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=144130 $D=1
M1347 936 933 1059 9 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=134870 $D=1
M1348 937 934 1060 9 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=139500 $D=1
M1349 938 935 1061 9 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=144130 $D=1
M1350 166 1 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=136120 $D=0
M1351 167 1 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=140750 $D=0
M1352 168 1 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=145380 $D=0
M1353 169 1 2 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=136120 $D=0
M1354 170 1 3 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=140750 $D=0
M1355 171 1 4 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=145380 $D=0
M1356 9 166 169 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=136120 $D=0
M1357 9 167 170 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=140750 $D=0
M1358 9 168 171 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=145380 $D=0
M1359 172 1 2 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=136120 $D=0
M1360 173 1 3 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=140750 $D=0
M1361 174 1 4 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=145380 $D=0
M1362 2 166 172 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=136120 $D=0
M1363 3 167 173 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=140750 $D=0
M1364 4 168 174 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=145380 $D=0
M1365 175 1 2 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=136120 $D=0
M1366 176 1 3 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=140750 $D=0
M1367 177 1 4 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=145380 $D=0
M1368 2 166 175 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=136120 $D=0
M1369 3 167 176 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=140750 $D=0
M1370 4 168 177 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=145380 $D=0
M1371 181 5 175 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=136120 $D=0
M1372 182 5 176 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=140750 $D=0
M1373 183 5 177 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=145380 $D=0
M1374 178 5 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=136120 $D=0
M1375 179 5 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=140750 $D=0
M1376 180 5 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=145380 $D=0
M1377 184 5 172 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=136120 $D=0
M1378 185 5 173 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=140750 $D=0
M1379 186 5 174 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=145380 $D=0
M1380 169 178 184 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=136120 $D=0
M1381 170 179 185 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=140750 $D=0
M1382 171 180 186 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=145380 $D=0
M1383 187 6 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=136120 $D=0
M1384 188 6 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=140750 $D=0
M1385 189 6 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=145380 $D=0
M1386 190 6 184 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=136120 $D=0
M1387 191 6 185 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=140750 $D=0
M1388 192 6 186 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=145380 $D=0
M1389 181 187 190 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=136120 $D=0
M1390 182 188 191 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=140750 $D=0
M1391 183 189 192 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=145380 $D=0
M1392 193 8 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=136120 $D=0
M1393 194 8 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=140750 $D=0
M1394 195 8 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=145380 $D=0
M1395 196 8 9 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=136120 $D=0
M1396 197 8 9 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=140750 $D=0
M1397 198 8 10 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=145380 $D=0
M1398 11 193 196 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=136120 $D=0
M1399 12 194 197 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=140750 $D=0
M1400 13 195 198 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=145380 $D=0
M1401 199 8 14 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=136120 $D=0
M1402 200 8 15 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=140750 $D=0
M1403 201 8 16 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=145380 $D=0
M1404 202 193 199 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=136120 $D=0
M1405 203 194 200 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=140750 $D=0
M1406 204 195 201 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=145380 $D=0
M1407 208 8 205 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=136120 $D=0
M1408 209 8 206 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=140750 $D=0
M1409 210 8 207 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=145380 $D=0
M1410 190 193 208 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=136120 $D=0
M1411 191 194 209 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=140750 $D=0
M1412 192 195 210 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=145380 $D=0
M1413 214 17 208 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=136120 $D=0
M1414 215 17 209 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=140750 $D=0
M1415 216 17 210 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=145380 $D=0
M1416 211 17 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=136120 $D=0
M1417 212 17 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=140750 $D=0
M1418 213 17 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=145380 $D=0
M1419 217 17 199 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=136120 $D=0
M1420 218 17 200 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=140750 $D=0
M1421 219 17 201 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=145380 $D=0
M1422 196 211 217 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=136120 $D=0
M1423 197 212 218 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=140750 $D=0
M1424 198 213 219 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=145380 $D=0
M1425 220 18 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=136120 $D=0
M1426 221 18 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=140750 $D=0
M1427 222 18 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=145380 $D=0
M1428 223 18 217 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=136120 $D=0
M1429 224 18 218 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=140750 $D=0
M1430 225 18 219 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=145380 $D=0
M1431 214 220 223 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=136120 $D=0
M1432 215 221 224 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=140750 $D=0
M1433 216 222 225 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=145380 $D=0
M1434 7 19 226 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=136120 $D=0
M1435 7 19 227 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=140750 $D=0
M1436 7 19 228 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=145380 $D=0
M1437 229 20 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=136120 $D=0
M1438 230 20 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=140750 $D=0
M1439 231 20 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=145380 $D=0
M1440 232 226 223 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=136120 $D=0
M1441 233 227 224 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=140750 $D=0
M1442 234 228 225 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=145380 $D=0
M1443 7 232 939 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=136120 $D=0
M1444 7 233 940 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=140750 $D=0
M1445 7 234 941 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=145380 $D=0
M1446 235 939 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=136120 $D=0
M1447 236 940 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=140750 $D=0
M1448 237 941 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=145380 $D=0
M1449 232 19 235 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=136120 $D=0
M1450 233 19 236 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=140750 $D=0
M1451 234 19 237 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=145380 $D=0
M1452 235 229 238 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=136120 $D=0
M1453 236 230 239 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=140750 $D=0
M1454 237 231 240 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=145380 $D=0
M1455 244 241 235 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=136120 $D=0
M1456 245 242 236 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=140750 $D=0
M1457 246 243 237 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=145380 $D=0
M1458 241 21 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=136120 $D=0
M1459 242 21 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=140750 $D=0
M1460 243 21 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=145380 $D=0
M1461 7 22 247 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=136120 $D=0
M1462 7 22 248 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=140750 $D=0
M1463 7 22 249 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=145380 $D=0
M1464 250 23 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=136120 $D=0
M1465 251 23 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=140750 $D=0
M1466 252 23 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=145380 $D=0
M1467 253 247 223 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=136120 $D=0
M1468 254 248 224 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=140750 $D=0
M1469 255 249 225 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=145380 $D=0
M1470 7 253 942 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=136120 $D=0
M1471 7 254 943 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=140750 $D=0
M1472 7 255 944 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=145380 $D=0
M1473 256 942 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=136120 $D=0
M1474 257 943 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=140750 $D=0
M1475 258 944 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=145380 $D=0
M1476 253 22 256 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=136120 $D=0
M1477 254 22 257 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=140750 $D=0
M1478 255 22 258 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=145380 $D=0
M1479 256 250 238 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=136120 $D=0
M1480 257 251 239 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=140750 $D=0
M1481 258 252 240 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=145380 $D=0
M1482 244 259 256 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=136120 $D=0
M1483 245 260 257 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=140750 $D=0
M1484 246 261 258 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=145380 $D=0
M1485 259 24 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=136120 $D=0
M1486 260 24 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=140750 $D=0
M1487 261 24 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=145380 $D=0
M1488 7 25 262 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=136120 $D=0
M1489 7 25 263 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=140750 $D=0
M1490 7 25 264 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=145380 $D=0
M1491 265 26 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=136120 $D=0
M1492 266 26 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=140750 $D=0
M1493 267 26 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=145380 $D=0
M1494 268 262 223 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=136120 $D=0
M1495 269 263 224 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=140750 $D=0
M1496 270 264 225 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=145380 $D=0
M1497 7 268 945 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=136120 $D=0
M1498 7 269 946 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=140750 $D=0
M1499 7 270 947 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=145380 $D=0
M1500 271 945 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=136120 $D=0
M1501 272 946 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=140750 $D=0
M1502 273 947 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=145380 $D=0
M1503 268 25 271 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=136120 $D=0
M1504 269 25 272 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=140750 $D=0
M1505 270 25 273 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=145380 $D=0
M1506 271 265 238 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=136120 $D=0
M1507 272 266 239 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=140750 $D=0
M1508 273 267 240 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=145380 $D=0
M1509 244 274 271 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=136120 $D=0
M1510 245 275 272 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=140750 $D=0
M1511 246 276 273 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=145380 $D=0
M1512 274 27 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=136120 $D=0
M1513 275 27 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=140750 $D=0
M1514 276 27 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=145380 $D=0
M1515 7 28 277 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=136120 $D=0
M1516 7 28 278 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=140750 $D=0
M1517 7 28 279 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=145380 $D=0
M1518 280 29 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=136120 $D=0
M1519 281 29 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=140750 $D=0
M1520 282 29 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=145380 $D=0
M1521 283 277 223 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=136120 $D=0
M1522 284 278 224 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=140750 $D=0
M1523 285 279 225 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=145380 $D=0
M1524 7 283 948 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=136120 $D=0
M1525 7 284 949 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=140750 $D=0
M1526 7 285 950 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=145380 $D=0
M1527 286 948 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=136120 $D=0
M1528 287 949 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=140750 $D=0
M1529 288 950 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=145380 $D=0
M1530 283 28 286 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=136120 $D=0
M1531 284 28 287 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=140750 $D=0
M1532 285 28 288 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=145380 $D=0
M1533 286 280 238 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=136120 $D=0
M1534 287 281 239 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=140750 $D=0
M1535 288 282 240 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=145380 $D=0
M1536 244 289 286 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=136120 $D=0
M1537 245 290 287 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=140750 $D=0
M1538 246 291 288 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=145380 $D=0
M1539 289 30 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=136120 $D=0
M1540 290 30 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=140750 $D=0
M1541 291 30 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=145380 $D=0
M1542 7 31 292 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=136120 $D=0
M1543 7 31 293 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=140750 $D=0
M1544 7 31 294 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=145380 $D=0
M1545 295 32 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=136120 $D=0
M1546 296 32 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=140750 $D=0
M1547 297 32 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=145380 $D=0
M1548 298 292 223 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=136120 $D=0
M1549 299 293 224 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=140750 $D=0
M1550 300 294 225 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=145380 $D=0
M1551 7 298 951 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=136120 $D=0
M1552 7 299 952 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=140750 $D=0
M1553 7 300 953 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=145380 $D=0
M1554 301 951 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=136120 $D=0
M1555 302 952 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=140750 $D=0
M1556 303 953 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=145380 $D=0
M1557 298 31 301 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=136120 $D=0
M1558 299 31 302 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=140750 $D=0
M1559 300 31 303 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=145380 $D=0
M1560 301 295 238 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=136120 $D=0
M1561 302 296 239 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=140750 $D=0
M1562 303 297 240 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=145380 $D=0
M1563 244 304 301 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=136120 $D=0
M1564 245 305 302 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=140750 $D=0
M1565 246 306 303 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=145380 $D=0
M1566 304 33 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=136120 $D=0
M1567 305 33 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=140750 $D=0
M1568 306 33 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=145380 $D=0
M1569 7 34 307 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=136120 $D=0
M1570 7 34 308 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=140750 $D=0
M1571 7 34 309 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=145380 $D=0
M1572 310 35 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=136120 $D=0
M1573 311 35 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=140750 $D=0
M1574 312 35 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=145380 $D=0
M1575 313 307 223 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=136120 $D=0
M1576 314 308 224 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=140750 $D=0
M1577 315 309 225 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=145380 $D=0
M1578 7 313 954 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=136120 $D=0
M1579 7 314 955 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=140750 $D=0
M1580 7 315 956 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=145380 $D=0
M1581 316 954 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=136120 $D=0
M1582 317 955 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=140750 $D=0
M1583 318 956 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=145380 $D=0
M1584 313 34 316 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=136120 $D=0
M1585 314 34 317 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=140750 $D=0
M1586 315 34 318 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=145380 $D=0
M1587 316 310 238 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=136120 $D=0
M1588 317 311 239 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=140750 $D=0
M1589 318 312 240 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=145380 $D=0
M1590 244 319 316 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=136120 $D=0
M1591 245 320 317 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=140750 $D=0
M1592 246 321 318 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=145380 $D=0
M1593 319 36 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=136120 $D=0
M1594 320 36 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=140750 $D=0
M1595 321 36 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=145380 $D=0
M1596 7 37 322 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=136120 $D=0
M1597 7 37 323 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=140750 $D=0
M1598 7 37 324 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=145380 $D=0
M1599 325 38 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=136120 $D=0
M1600 326 38 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=140750 $D=0
M1601 327 38 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=145380 $D=0
M1602 328 322 223 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=136120 $D=0
M1603 329 323 224 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=140750 $D=0
M1604 330 324 225 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=145380 $D=0
M1605 7 328 957 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=136120 $D=0
M1606 7 329 958 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=140750 $D=0
M1607 7 330 959 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=145380 $D=0
M1608 331 957 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=136120 $D=0
M1609 332 958 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=140750 $D=0
M1610 333 959 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=145380 $D=0
M1611 328 37 331 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=136120 $D=0
M1612 329 37 332 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=140750 $D=0
M1613 330 37 333 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=145380 $D=0
M1614 331 325 238 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=136120 $D=0
M1615 332 326 239 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=140750 $D=0
M1616 333 327 240 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=145380 $D=0
M1617 244 334 331 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=136120 $D=0
M1618 245 335 332 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=140750 $D=0
M1619 246 336 333 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=145380 $D=0
M1620 334 39 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=136120 $D=0
M1621 335 39 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=140750 $D=0
M1622 336 39 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=145380 $D=0
M1623 7 40 337 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=136120 $D=0
M1624 7 40 338 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=140750 $D=0
M1625 7 40 339 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=145380 $D=0
M1626 340 41 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=136120 $D=0
M1627 341 41 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=140750 $D=0
M1628 342 41 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=145380 $D=0
M1629 343 337 223 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=136120 $D=0
M1630 344 338 224 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=140750 $D=0
M1631 345 339 225 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=145380 $D=0
M1632 7 343 960 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=136120 $D=0
M1633 7 344 961 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=140750 $D=0
M1634 7 345 962 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=145380 $D=0
M1635 346 960 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=136120 $D=0
M1636 347 961 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=140750 $D=0
M1637 348 962 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=145380 $D=0
M1638 343 40 346 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=136120 $D=0
M1639 344 40 347 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=140750 $D=0
M1640 345 40 348 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=145380 $D=0
M1641 346 340 238 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=136120 $D=0
M1642 347 341 239 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=140750 $D=0
M1643 348 342 240 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=145380 $D=0
M1644 244 349 346 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=136120 $D=0
M1645 245 350 347 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=140750 $D=0
M1646 246 351 348 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=145380 $D=0
M1647 349 42 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=136120 $D=0
M1648 350 42 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=140750 $D=0
M1649 351 42 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=145380 $D=0
M1650 7 43 352 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=136120 $D=0
M1651 7 43 353 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=140750 $D=0
M1652 7 43 354 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=145380 $D=0
M1653 355 44 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=136120 $D=0
M1654 356 44 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=140750 $D=0
M1655 357 44 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=145380 $D=0
M1656 358 352 223 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=136120 $D=0
M1657 359 353 224 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=140750 $D=0
M1658 360 354 225 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=145380 $D=0
M1659 7 358 963 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=136120 $D=0
M1660 7 359 964 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=140750 $D=0
M1661 7 360 965 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=145380 $D=0
M1662 361 963 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=136120 $D=0
M1663 362 964 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=140750 $D=0
M1664 363 965 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=145380 $D=0
M1665 358 43 361 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=136120 $D=0
M1666 359 43 362 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=140750 $D=0
M1667 360 43 363 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=145380 $D=0
M1668 361 355 238 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=136120 $D=0
M1669 362 356 239 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=140750 $D=0
M1670 363 357 240 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=145380 $D=0
M1671 244 364 361 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=136120 $D=0
M1672 245 365 362 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=140750 $D=0
M1673 246 366 363 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=145380 $D=0
M1674 364 45 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=136120 $D=0
M1675 365 45 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=140750 $D=0
M1676 366 45 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=145380 $D=0
M1677 7 46 367 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=136120 $D=0
M1678 7 46 368 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=140750 $D=0
M1679 7 46 369 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=145380 $D=0
M1680 370 47 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=136120 $D=0
M1681 371 47 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=140750 $D=0
M1682 372 47 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=145380 $D=0
M1683 373 367 223 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=136120 $D=0
M1684 374 368 224 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=140750 $D=0
M1685 375 369 225 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=145380 $D=0
M1686 7 373 966 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=136120 $D=0
M1687 7 374 967 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=140750 $D=0
M1688 7 375 968 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=145380 $D=0
M1689 376 966 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=136120 $D=0
M1690 377 967 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=140750 $D=0
M1691 378 968 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=145380 $D=0
M1692 373 46 376 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=136120 $D=0
M1693 374 46 377 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=140750 $D=0
M1694 375 46 378 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=145380 $D=0
M1695 376 370 238 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=136120 $D=0
M1696 377 371 239 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=140750 $D=0
M1697 378 372 240 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=145380 $D=0
M1698 244 379 376 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=136120 $D=0
M1699 245 380 377 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=140750 $D=0
M1700 246 381 378 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=145380 $D=0
M1701 379 48 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=136120 $D=0
M1702 380 48 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=140750 $D=0
M1703 381 48 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=145380 $D=0
M1704 7 49 382 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=136120 $D=0
M1705 7 49 383 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=140750 $D=0
M1706 7 49 384 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=145380 $D=0
M1707 385 50 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=136120 $D=0
M1708 386 50 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=140750 $D=0
M1709 387 50 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=145380 $D=0
M1710 388 382 223 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=136120 $D=0
M1711 389 383 224 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=140750 $D=0
M1712 390 384 225 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=145380 $D=0
M1713 7 388 969 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=136120 $D=0
M1714 7 389 970 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=140750 $D=0
M1715 7 390 971 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=145380 $D=0
M1716 391 969 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=136120 $D=0
M1717 392 970 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=140750 $D=0
M1718 393 971 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=145380 $D=0
M1719 388 49 391 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=136120 $D=0
M1720 389 49 392 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=140750 $D=0
M1721 390 49 393 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=145380 $D=0
M1722 391 385 238 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=136120 $D=0
M1723 392 386 239 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=140750 $D=0
M1724 393 387 240 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=145380 $D=0
M1725 244 394 391 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=136120 $D=0
M1726 245 395 392 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=140750 $D=0
M1727 246 396 393 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=145380 $D=0
M1728 394 51 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=136120 $D=0
M1729 395 51 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=140750 $D=0
M1730 396 51 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=145380 $D=0
M1731 7 52 397 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=136120 $D=0
M1732 7 52 398 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=140750 $D=0
M1733 7 52 399 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=145380 $D=0
M1734 400 53 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=136120 $D=0
M1735 401 53 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=140750 $D=0
M1736 402 53 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=145380 $D=0
M1737 403 397 223 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=136120 $D=0
M1738 404 398 224 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=140750 $D=0
M1739 405 399 225 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=145380 $D=0
M1740 7 403 972 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=136120 $D=0
M1741 7 404 973 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=140750 $D=0
M1742 7 405 974 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=145380 $D=0
M1743 406 972 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=136120 $D=0
M1744 407 973 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=140750 $D=0
M1745 408 974 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=145380 $D=0
M1746 403 52 406 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=136120 $D=0
M1747 404 52 407 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=140750 $D=0
M1748 405 52 408 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=145380 $D=0
M1749 406 400 238 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=136120 $D=0
M1750 407 401 239 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=140750 $D=0
M1751 408 402 240 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=145380 $D=0
M1752 244 409 406 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=136120 $D=0
M1753 245 410 407 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=140750 $D=0
M1754 246 411 408 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=145380 $D=0
M1755 409 54 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=136120 $D=0
M1756 410 54 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=140750 $D=0
M1757 411 54 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=145380 $D=0
M1758 7 55 412 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=136120 $D=0
M1759 7 55 413 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=140750 $D=0
M1760 7 55 414 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=145380 $D=0
M1761 415 56 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=136120 $D=0
M1762 416 56 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=140750 $D=0
M1763 417 56 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=145380 $D=0
M1764 418 412 223 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=136120 $D=0
M1765 419 413 224 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=140750 $D=0
M1766 420 414 225 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=145380 $D=0
M1767 7 418 975 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=136120 $D=0
M1768 7 419 976 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=140750 $D=0
M1769 7 420 977 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=145380 $D=0
M1770 421 975 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=136120 $D=0
M1771 422 976 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=140750 $D=0
M1772 423 977 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=145380 $D=0
M1773 418 55 421 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=136120 $D=0
M1774 419 55 422 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=140750 $D=0
M1775 420 55 423 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=145380 $D=0
M1776 421 415 238 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=136120 $D=0
M1777 422 416 239 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=140750 $D=0
M1778 423 417 240 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=145380 $D=0
M1779 244 424 421 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=136120 $D=0
M1780 245 425 422 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=140750 $D=0
M1781 246 426 423 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=145380 $D=0
M1782 424 57 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=136120 $D=0
M1783 425 57 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=140750 $D=0
M1784 426 57 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=145380 $D=0
M1785 7 58 427 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=136120 $D=0
M1786 7 58 428 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=140750 $D=0
M1787 7 58 429 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=145380 $D=0
M1788 430 59 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=136120 $D=0
M1789 431 59 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=140750 $D=0
M1790 432 59 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=145380 $D=0
M1791 433 427 223 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=136120 $D=0
M1792 434 428 224 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=140750 $D=0
M1793 435 429 225 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=145380 $D=0
M1794 7 433 978 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=136120 $D=0
M1795 7 434 979 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=140750 $D=0
M1796 7 435 980 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=145380 $D=0
M1797 436 978 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=136120 $D=0
M1798 437 979 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=140750 $D=0
M1799 438 980 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=145380 $D=0
M1800 433 58 436 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=136120 $D=0
M1801 434 58 437 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=140750 $D=0
M1802 435 58 438 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=145380 $D=0
M1803 436 430 238 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=136120 $D=0
M1804 437 431 239 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=140750 $D=0
M1805 438 432 240 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=145380 $D=0
M1806 244 439 436 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=136120 $D=0
M1807 245 440 437 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=140750 $D=0
M1808 246 441 438 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=145380 $D=0
M1809 439 60 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=136120 $D=0
M1810 440 60 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=140750 $D=0
M1811 441 60 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=145380 $D=0
M1812 7 61 442 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=136120 $D=0
M1813 7 61 443 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=140750 $D=0
M1814 7 61 444 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=145380 $D=0
M1815 445 62 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=136120 $D=0
M1816 446 62 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=140750 $D=0
M1817 447 62 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=145380 $D=0
M1818 448 442 223 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=136120 $D=0
M1819 449 443 224 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=140750 $D=0
M1820 450 444 225 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=145380 $D=0
M1821 7 448 981 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=136120 $D=0
M1822 7 449 982 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=140750 $D=0
M1823 7 450 983 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=145380 $D=0
M1824 451 981 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=136120 $D=0
M1825 452 982 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=140750 $D=0
M1826 453 983 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=145380 $D=0
M1827 448 61 451 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=136120 $D=0
M1828 449 61 452 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=140750 $D=0
M1829 450 61 453 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=145380 $D=0
M1830 451 445 238 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=136120 $D=0
M1831 452 446 239 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=140750 $D=0
M1832 453 447 240 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=145380 $D=0
M1833 244 454 451 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=136120 $D=0
M1834 245 455 452 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=140750 $D=0
M1835 246 456 453 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=145380 $D=0
M1836 454 63 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=136120 $D=0
M1837 455 63 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=140750 $D=0
M1838 456 63 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=145380 $D=0
M1839 7 64 457 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=136120 $D=0
M1840 7 64 458 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=140750 $D=0
M1841 7 64 459 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=145380 $D=0
M1842 460 65 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=136120 $D=0
M1843 461 65 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=140750 $D=0
M1844 462 65 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=145380 $D=0
M1845 463 457 223 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=136120 $D=0
M1846 464 458 224 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=140750 $D=0
M1847 465 459 225 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=145380 $D=0
M1848 7 463 984 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=136120 $D=0
M1849 7 464 985 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=140750 $D=0
M1850 7 465 986 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=145380 $D=0
M1851 466 984 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=136120 $D=0
M1852 467 985 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=140750 $D=0
M1853 468 986 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=145380 $D=0
M1854 463 64 466 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=136120 $D=0
M1855 464 64 467 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=140750 $D=0
M1856 465 64 468 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=145380 $D=0
M1857 466 460 238 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=136120 $D=0
M1858 467 461 239 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=140750 $D=0
M1859 468 462 240 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=145380 $D=0
M1860 244 469 466 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=136120 $D=0
M1861 245 470 467 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=140750 $D=0
M1862 246 471 468 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=145380 $D=0
M1863 469 66 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=136120 $D=0
M1864 470 66 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=140750 $D=0
M1865 471 66 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=145380 $D=0
M1866 7 67 472 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=136120 $D=0
M1867 7 67 473 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=140750 $D=0
M1868 7 67 474 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=145380 $D=0
M1869 475 68 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=136120 $D=0
M1870 476 68 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=140750 $D=0
M1871 477 68 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=145380 $D=0
M1872 478 472 223 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=136120 $D=0
M1873 479 473 224 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=140750 $D=0
M1874 480 474 225 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=145380 $D=0
M1875 7 478 987 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=136120 $D=0
M1876 7 479 988 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=140750 $D=0
M1877 7 480 989 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=145380 $D=0
M1878 481 987 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=136120 $D=0
M1879 482 988 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=140750 $D=0
M1880 483 989 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=145380 $D=0
M1881 478 67 481 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=136120 $D=0
M1882 479 67 482 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=140750 $D=0
M1883 480 67 483 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=145380 $D=0
M1884 481 475 238 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=136120 $D=0
M1885 482 476 239 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=140750 $D=0
M1886 483 477 240 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=145380 $D=0
M1887 244 484 481 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=136120 $D=0
M1888 245 485 482 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=140750 $D=0
M1889 246 486 483 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=145380 $D=0
M1890 484 69 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=136120 $D=0
M1891 485 69 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=140750 $D=0
M1892 486 69 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=145380 $D=0
M1893 7 70 487 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=136120 $D=0
M1894 7 70 488 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=140750 $D=0
M1895 7 70 489 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=145380 $D=0
M1896 490 71 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=136120 $D=0
M1897 491 71 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=140750 $D=0
M1898 492 71 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=145380 $D=0
M1899 493 487 223 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=136120 $D=0
M1900 494 488 224 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=140750 $D=0
M1901 495 489 225 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=145380 $D=0
M1902 7 493 990 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=136120 $D=0
M1903 7 494 991 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=140750 $D=0
M1904 7 495 992 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=145380 $D=0
M1905 496 990 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=136120 $D=0
M1906 497 991 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=140750 $D=0
M1907 498 992 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=145380 $D=0
M1908 493 70 496 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=136120 $D=0
M1909 494 70 497 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=140750 $D=0
M1910 495 70 498 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=145380 $D=0
M1911 496 490 238 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=136120 $D=0
M1912 497 491 239 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=140750 $D=0
M1913 498 492 240 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=145380 $D=0
M1914 244 499 496 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=136120 $D=0
M1915 245 500 497 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=140750 $D=0
M1916 246 501 498 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=145380 $D=0
M1917 499 72 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=136120 $D=0
M1918 500 72 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=140750 $D=0
M1919 501 72 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=145380 $D=0
M1920 7 73 502 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=136120 $D=0
M1921 7 73 503 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=140750 $D=0
M1922 7 73 504 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=145380 $D=0
M1923 505 74 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=136120 $D=0
M1924 506 74 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=140750 $D=0
M1925 507 74 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=145380 $D=0
M1926 508 502 223 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=136120 $D=0
M1927 509 503 224 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=140750 $D=0
M1928 510 504 225 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=145380 $D=0
M1929 7 508 993 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=136120 $D=0
M1930 7 509 994 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=140750 $D=0
M1931 7 510 995 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=145380 $D=0
M1932 511 993 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=136120 $D=0
M1933 512 994 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=140750 $D=0
M1934 513 995 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=145380 $D=0
M1935 508 73 511 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=136120 $D=0
M1936 509 73 512 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=140750 $D=0
M1937 510 73 513 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=145380 $D=0
M1938 511 505 238 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=136120 $D=0
M1939 512 506 239 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=140750 $D=0
M1940 513 507 240 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=145380 $D=0
M1941 244 514 511 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=136120 $D=0
M1942 245 515 512 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=140750 $D=0
M1943 246 516 513 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=145380 $D=0
M1944 514 75 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=136120 $D=0
M1945 515 75 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=140750 $D=0
M1946 516 75 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=145380 $D=0
M1947 7 76 517 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=136120 $D=0
M1948 7 76 518 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=140750 $D=0
M1949 7 76 519 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=145380 $D=0
M1950 520 77 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=136120 $D=0
M1951 521 77 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=140750 $D=0
M1952 522 77 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=145380 $D=0
M1953 523 517 223 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=136120 $D=0
M1954 524 518 224 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=140750 $D=0
M1955 525 519 225 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=145380 $D=0
M1956 7 523 996 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=136120 $D=0
M1957 7 524 997 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=140750 $D=0
M1958 7 525 998 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=145380 $D=0
M1959 526 996 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=136120 $D=0
M1960 527 997 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=140750 $D=0
M1961 528 998 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=145380 $D=0
M1962 523 76 526 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=136120 $D=0
M1963 524 76 527 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=140750 $D=0
M1964 525 76 528 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=145380 $D=0
M1965 526 520 238 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=136120 $D=0
M1966 527 521 239 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=140750 $D=0
M1967 528 522 240 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=145380 $D=0
M1968 244 529 526 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=136120 $D=0
M1969 245 530 527 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=140750 $D=0
M1970 246 531 528 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=145380 $D=0
M1971 529 78 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=136120 $D=0
M1972 530 78 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=140750 $D=0
M1973 531 78 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=145380 $D=0
M1974 7 79 532 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=136120 $D=0
M1975 7 79 533 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=140750 $D=0
M1976 7 79 534 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=145380 $D=0
M1977 535 80 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=136120 $D=0
M1978 536 80 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=140750 $D=0
M1979 537 80 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=145380 $D=0
M1980 538 532 223 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=136120 $D=0
M1981 539 533 224 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=140750 $D=0
M1982 540 534 225 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=145380 $D=0
M1983 7 538 999 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=136120 $D=0
M1984 7 539 1000 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=140750 $D=0
M1985 7 540 1001 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=145380 $D=0
M1986 541 999 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=136120 $D=0
M1987 542 1000 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=140750 $D=0
M1988 543 1001 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=145380 $D=0
M1989 538 79 541 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=136120 $D=0
M1990 539 79 542 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=140750 $D=0
M1991 540 79 543 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=145380 $D=0
M1992 541 535 238 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=136120 $D=0
M1993 542 536 239 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=140750 $D=0
M1994 543 537 240 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=145380 $D=0
M1995 244 544 541 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=136120 $D=0
M1996 245 545 542 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=140750 $D=0
M1997 246 546 543 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=145380 $D=0
M1998 544 81 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=136120 $D=0
M1999 545 81 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=140750 $D=0
M2000 546 81 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=145380 $D=0
M2001 7 82 547 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=136120 $D=0
M2002 7 82 548 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=140750 $D=0
M2003 7 82 549 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=145380 $D=0
M2004 550 83 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=136120 $D=0
M2005 551 83 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=140750 $D=0
M2006 552 83 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=145380 $D=0
M2007 553 547 223 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=136120 $D=0
M2008 554 548 224 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=140750 $D=0
M2009 555 549 225 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=145380 $D=0
M2010 7 553 1002 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=136120 $D=0
M2011 7 554 1003 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=140750 $D=0
M2012 7 555 1004 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=145380 $D=0
M2013 556 1002 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=136120 $D=0
M2014 557 1003 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=140750 $D=0
M2015 558 1004 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=145380 $D=0
M2016 553 82 556 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=136120 $D=0
M2017 554 82 557 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=140750 $D=0
M2018 555 82 558 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=145380 $D=0
M2019 556 550 238 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=136120 $D=0
M2020 557 551 239 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=140750 $D=0
M2021 558 552 240 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=145380 $D=0
M2022 244 559 556 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=136120 $D=0
M2023 245 560 557 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=140750 $D=0
M2024 246 561 558 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=145380 $D=0
M2025 559 84 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=136120 $D=0
M2026 560 84 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=140750 $D=0
M2027 561 84 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=145380 $D=0
M2028 7 85 562 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=136120 $D=0
M2029 7 85 563 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=140750 $D=0
M2030 7 85 564 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=145380 $D=0
M2031 565 86 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=136120 $D=0
M2032 566 86 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=140750 $D=0
M2033 567 86 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=145380 $D=0
M2034 568 562 223 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=136120 $D=0
M2035 569 563 224 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=140750 $D=0
M2036 570 564 225 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=145380 $D=0
M2037 7 568 1005 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=136120 $D=0
M2038 7 569 1006 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=140750 $D=0
M2039 7 570 1007 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=145380 $D=0
M2040 571 1005 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=136120 $D=0
M2041 572 1006 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=140750 $D=0
M2042 573 1007 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=145380 $D=0
M2043 568 85 571 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=136120 $D=0
M2044 569 85 572 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=140750 $D=0
M2045 570 85 573 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=145380 $D=0
M2046 571 565 238 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=136120 $D=0
M2047 572 566 239 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=140750 $D=0
M2048 573 567 240 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=145380 $D=0
M2049 244 574 571 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=136120 $D=0
M2050 245 575 572 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=140750 $D=0
M2051 246 576 573 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=145380 $D=0
M2052 574 87 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=136120 $D=0
M2053 575 87 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=140750 $D=0
M2054 576 87 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=145380 $D=0
M2055 7 88 577 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=136120 $D=0
M2056 7 88 578 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=140750 $D=0
M2057 7 88 579 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=145380 $D=0
M2058 580 89 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=136120 $D=0
M2059 581 89 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=140750 $D=0
M2060 582 89 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=145380 $D=0
M2061 583 577 223 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=136120 $D=0
M2062 584 578 224 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=140750 $D=0
M2063 585 579 225 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=145380 $D=0
M2064 7 583 1008 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=136120 $D=0
M2065 7 584 1009 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=140750 $D=0
M2066 7 585 1010 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=145380 $D=0
M2067 586 1008 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=136120 $D=0
M2068 587 1009 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=140750 $D=0
M2069 588 1010 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=145380 $D=0
M2070 583 88 586 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=136120 $D=0
M2071 584 88 587 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=140750 $D=0
M2072 585 88 588 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=145380 $D=0
M2073 586 580 238 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=136120 $D=0
M2074 587 581 239 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=140750 $D=0
M2075 588 582 240 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=145380 $D=0
M2076 244 589 586 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=136120 $D=0
M2077 245 590 587 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=140750 $D=0
M2078 246 591 588 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=145380 $D=0
M2079 589 90 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=136120 $D=0
M2080 590 90 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=140750 $D=0
M2081 591 90 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=145380 $D=0
M2082 7 91 592 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=136120 $D=0
M2083 7 91 593 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=140750 $D=0
M2084 7 91 594 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=145380 $D=0
M2085 595 92 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=136120 $D=0
M2086 596 92 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=140750 $D=0
M2087 597 92 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=145380 $D=0
M2088 598 592 223 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=136120 $D=0
M2089 599 593 224 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=140750 $D=0
M2090 600 594 225 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=145380 $D=0
M2091 7 598 1011 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=136120 $D=0
M2092 7 599 1012 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=140750 $D=0
M2093 7 600 1013 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=145380 $D=0
M2094 601 1011 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=136120 $D=0
M2095 602 1012 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=140750 $D=0
M2096 603 1013 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=145380 $D=0
M2097 598 91 601 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=136120 $D=0
M2098 599 91 602 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=140750 $D=0
M2099 600 91 603 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=145380 $D=0
M2100 601 595 238 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=136120 $D=0
M2101 602 596 239 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=140750 $D=0
M2102 603 597 240 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=145380 $D=0
M2103 244 604 601 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=136120 $D=0
M2104 245 605 602 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=140750 $D=0
M2105 246 606 603 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=145380 $D=0
M2106 604 93 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=136120 $D=0
M2107 605 93 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=140750 $D=0
M2108 606 93 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=145380 $D=0
M2109 7 94 607 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=136120 $D=0
M2110 7 94 608 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=140750 $D=0
M2111 7 94 609 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=145380 $D=0
M2112 610 95 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=136120 $D=0
M2113 611 95 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=140750 $D=0
M2114 612 95 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=145380 $D=0
M2115 613 607 223 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=136120 $D=0
M2116 614 608 224 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=140750 $D=0
M2117 615 609 225 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=145380 $D=0
M2118 7 613 1014 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=136120 $D=0
M2119 7 614 1015 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=140750 $D=0
M2120 7 615 1016 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=145380 $D=0
M2121 616 1014 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=136120 $D=0
M2122 617 1015 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=140750 $D=0
M2123 618 1016 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=145380 $D=0
M2124 613 94 616 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=136120 $D=0
M2125 614 94 617 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=140750 $D=0
M2126 615 94 618 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=145380 $D=0
M2127 616 610 238 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=136120 $D=0
M2128 617 611 239 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=140750 $D=0
M2129 618 612 240 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=145380 $D=0
M2130 244 619 616 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=136120 $D=0
M2131 245 620 617 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=140750 $D=0
M2132 246 621 618 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=145380 $D=0
M2133 619 96 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=136120 $D=0
M2134 620 96 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=140750 $D=0
M2135 621 96 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=145380 $D=0
M2136 7 97 622 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=136120 $D=0
M2137 7 97 623 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=140750 $D=0
M2138 7 97 624 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=145380 $D=0
M2139 625 98 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=136120 $D=0
M2140 626 98 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=140750 $D=0
M2141 627 98 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=145380 $D=0
M2142 628 622 223 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=136120 $D=0
M2143 629 623 224 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=140750 $D=0
M2144 630 624 225 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=145380 $D=0
M2145 7 628 1017 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=136120 $D=0
M2146 7 629 1018 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=140750 $D=0
M2147 7 630 1019 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=145380 $D=0
M2148 631 1017 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=136120 $D=0
M2149 632 1018 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=140750 $D=0
M2150 633 1019 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=145380 $D=0
M2151 628 97 631 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=136120 $D=0
M2152 629 97 632 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=140750 $D=0
M2153 630 97 633 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=145380 $D=0
M2154 631 625 238 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=136120 $D=0
M2155 632 626 239 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=140750 $D=0
M2156 633 627 240 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=145380 $D=0
M2157 244 634 631 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=136120 $D=0
M2158 245 635 632 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=140750 $D=0
M2159 246 636 633 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=145380 $D=0
M2160 634 99 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=136120 $D=0
M2161 635 99 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=140750 $D=0
M2162 636 99 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=145380 $D=0
M2163 7 100 637 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=136120 $D=0
M2164 7 100 638 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=140750 $D=0
M2165 7 100 639 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=145380 $D=0
M2166 640 101 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=136120 $D=0
M2167 641 101 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=140750 $D=0
M2168 642 101 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=145380 $D=0
M2169 643 637 223 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=136120 $D=0
M2170 644 638 224 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=140750 $D=0
M2171 645 639 225 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=145380 $D=0
M2172 7 643 1020 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=136120 $D=0
M2173 7 644 1021 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=140750 $D=0
M2174 7 645 1022 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=145380 $D=0
M2175 646 1020 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=136120 $D=0
M2176 647 1021 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=140750 $D=0
M2177 648 1022 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=145380 $D=0
M2178 643 100 646 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=136120 $D=0
M2179 644 100 647 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=140750 $D=0
M2180 645 100 648 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=145380 $D=0
M2181 646 640 238 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=136120 $D=0
M2182 647 641 239 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=140750 $D=0
M2183 648 642 240 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=145380 $D=0
M2184 244 649 646 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=136120 $D=0
M2185 245 650 647 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=140750 $D=0
M2186 246 651 648 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=145380 $D=0
M2187 649 102 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=136120 $D=0
M2188 650 102 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=140750 $D=0
M2189 651 102 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=145380 $D=0
M2190 7 103 652 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=136120 $D=0
M2191 7 103 653 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=140750 $D=0
M2192 7 103 654 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=145380 $D=0
M2193 655 104 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=136120 $D=0
M2194 656 104 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=140750 $D=0
M2195 657 104 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=145380 $D=0
M2196 658 652 223 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=136120 $D=0
M2197 659 653 224 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=140750 $D=0
M2198 660 654 225 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=145380 $D=0
M2199 7 658 1023 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=136120 $D=0
M2200 7 659 1024 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=140750 $D=0
M2201 7 660 1025 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=145380 $D=0
M2202 661 1023 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=136120 $D=0
M2203 662 1024 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=140750 $D=0
M2204 663 1025 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=145380 $D=0
M2205 658 103 661 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=136120 $D=0
M2206 659 103 662 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=140750 $D=0
M2207 660 103 663 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=145380 $D=0
M2208 661 655 238 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=136120 $D=0
M2209 662 656 239 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=140750 $D=0
M2210 663 657 240 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=145380 $D=0
M2211 244 664 661 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=136120 $D=0
M2212 245 665 662 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=140750 $D=0
M2213 246 666 663 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=145380 $D=0
M2214 664 105 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=136120 $D=0
M2215 665 105 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=140750 $D=0
M2216 666 105 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=145380 $D=0
M2217 7 106 667 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=136120 $D=0
M2218 7 106 668 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=140750 $D=0
M2219 7 106 669 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=145380 $D=0
M2220 670 107 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=136120 $D=0
M2221 671 107 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=140750 $D=0
M2222 672 107 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=145380 $D=0
M2223 673 667 223 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=136120 $D=0
M2224 674 668 224 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=140750 $D=0
M2225 675 669 225 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=145380 $D=0
M2226 7 673 1026 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=136120 $D=0
M2227 7 674 1027 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=140750 $D=0
M2228 7 675 1028 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=145380 $D=0
M2229 676 1026 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=136120 $D=0
M2230 677 1027 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=140750 $D=0
M2231 678 1028 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=145380 $D=0
M2232 673 106 676 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=136120 $D=0
M2233 674 106 677 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=140750 $D=0
M2234 675 106 678 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=145380 $D=0
M2235 676 670 238 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=136120 $D=0
M2236 677 671 239 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=140750 $D=0
M2237 678 672 240 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=145380 $D=0
M2238 244 679 676 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=136120 $D=0
M2239 245 680 677 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=140750 $D=0
M2240 246 681 678 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=145380 $D=0
M2241 679 108 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=136120 $D=0
M2242 680 108 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=140750 $D=0
M2243 681 108 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=145380 $D=0
M2244 7 109 682 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=136120 $D=0
M2245 7 109 683 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=140750 $D=0
M2246 7 109 684 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=145380 $D=0
M2247 685 110 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=136120 $D=0
M2248 686 110 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=140750 $D=0
M2249 687 110 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=145380 $D=0
M2250 688 682 223 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=136120 $D=0
M2251 689 683 224 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=140750 $D=0
M2252 690 684 225 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=145380 $D=0
M2253 7 688 1029 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=136120 $D=0
M2254 7 689 1030 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=140750 $D=0
M2255 7 690 1031 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=145380 $D=0
M2256 691 1029 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=136120 $D=0
M2257 692 1030 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=140750 $D=0
M2258 693 1031 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=145380 $D=0
M2259 688 109 691 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=136120 $D=0
M2260 689 109 692 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=140750 $D=0
M2261 690 109 693 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=145380 $D=0
M2262 691 685 238 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=136120 $D=0
M2263 692 686 239 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=140750 $D=0
M2264 693 687 240 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=145380 $D=0
M2265 244 694 691 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=136120 $D=0
M2266 245 695 692 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=140750 $D=0
M2267 246 696 693 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=145380 $D=0
M2268 694 111 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=136120 $D=0
M2269 695 111 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=140750 $D=0
M2270 696 111 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=145380 $D=0
M2271 7 112 697 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=136120 $D=0
M2272 7 112 698 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=140750 $D=0
M2273 7 112 699 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=145380 $D=0
M2274 700 113 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=136120 $D=0
M2275 701 113 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=140750 $D=0
M2276 702 113 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=145380 $D=0
M2277 9 700 238 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=136120 $D=0
M2278 9 701 239 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=140750 $D=0
M2279 9 702 240 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=145380 $D=0
M2280 244 697 9 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=136120 $D=0
M2281 245 698 9 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=140750 $D=0
M2282 246 699 9 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=145380 $D=0
M2283 7 706 703 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=136120 $D=0
M2284 7 707 704 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=140750 $D=0
M2285 7 708 705 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=145380 $D=0
M2286 706 114 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=136120 $D=0
M2287 707 114 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=140750 $D=0
M2288 708 114 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=145380 $D=0
M2289 1032 238 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=136120 $D=0
M2290 1033 239 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=140750 $D=0
M2291 1034 240 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=145380 $D=0
M2292 709 706 1032 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=136120 $D=0
M2293 710 707 1033 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=140750 $D=0
M2294 711 708 1034 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=145380 $D=0
M2295 7 709 712 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=136120 $D=0
M2296 7 710 713 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=140750 $D=0
M2297 7 711 714 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=145380 $D=0
M2298 1035 712 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=136120 $D=0
M2299 1036 713 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=140750 $D=0
M2300 1037 714 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=145380 $D=0
M2301 709 703 1035 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=136120 $D=0
M2302 710 704 1036 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=140750 $D=0
M2303 711 705 1037 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=145380 $D=0
M2304 7 718 715 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=136120 $D=0
M2305 7 719 716 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=140750 $D=0
M2306 7 720 717 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=145380 $D=0
M2307 718 114 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=136120 $D=0
M2308 719 114 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=140750 $D=0
M2309 720 114 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=145380 $D=0
M2310 1038 244 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=136120 $D=0
M2311 1039 245 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=140750 $D=0
M2312 1040 246 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=145380 $D=0
M2313 721 718 1038 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=136120 $D=0
M2314 722 719 1039 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=140750 $D=0
M2315 723 720 1040 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=145380 $D=0
M2316 7 721 115 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=136120 $D=0
M2317 7 722 116 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=140750 $D=0
M2318 7 723 117 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=145380 $D=0
M2319 1041 115 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=136120 $D=0
M2320 1042 116 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=140750 $D=0
M2321 1043 117 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=145380 $D=0
M2322 721 715 1041 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=136120 $D=0
M2323 722 716 1042 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=140750 $D=0
M2324 723 717 1043 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=145380 $D=0
M2325 724 118 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=136120 $D=0
M2326 725 118 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=140750 $D=0
M2327 726 118 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=145380 $D=0
M2328 727 118 712 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=136120 $D=0
M2329 728 118 713 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=140750 $D=0
M2330 729 118 714 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=145380 $D=0
M2331 119 724 727 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=136120 $D=0
M2332 120 725 728 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=140750 $D=0
M2333 121 726 729 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=145380 $D=0
M2334 730 122 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=136120 $D=0
M2335 731 122 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=140750 $D=0
M2336 732 122 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=145380 $D=0
M2337 733 122 115 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=136120 $D=0
M2338 734 122 116 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=140750 $D=0
M2339 735 122 117 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=145380 $D=0
M2340 1044 730 733 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=136120 $D=0
M2341 1045 731 734 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=140750 $D=0
M2342 1046 732 735 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=145380 $D=0
M2343 7 115 1044 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=136120 $D=0
M2344 7 116 1045 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=140750 $D=0
M2345 7 117 1046 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=145380 $D=0
M2346 736 123 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=136120 $D=0
M2347 737 123 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=140750 $D=0
M2348 738 123 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=145380 $D=0
M2349 124 123 733 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=136120 $D=0
M2350 125 123 734 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=140750 $D=0
M2351 126 123 735 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=145380 $D=0
M2352 11 736 124 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=136120 $D=0
M2353 12 737 125 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=140750 $D=0
M2354 13 738 126 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=145380 $D=0
M2355 741 739 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=136120 $D=0
M2356 742 740 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=140750 $D=0
M2357 743 127 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=145380 $D=0
M2358 7 747 744 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=136120 $D=0
M2359 7 748 745 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=140750 $D=0
M2360 7 749 746 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=145380 $D=0
M2361 750 727 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=136120 $D=0
M2362 751 728 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=140750 $D=0
M2363 752 729 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=145380 $D=0
M2364 747 727 739 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=136120 $D=0
M2365 748 728 740 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=140750 $D=0
M2366 749 729 127 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=145380 $D=0
M2367 741 750 747 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=136120 $D=0
M2368 742 751 748 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=140750 $D=0
M2369 743 752 749 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=145380 $D=0
M2370 753 744 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=136120 $D=0
M2371 754 745 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=140750 $D=0
M2372 755 746 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=145380 $D=0
M2373 128 744 124 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=136120 $D=0
M2374 739 745 125 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=140750 $D=0
M2375 740 746 126 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=145380 $D=0
M2376 727 753 128 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=136120 $D=0
M2377 728 754 739 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=140750 $D=0
M2378 729 755 740 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=145380 $D=0
M2379 756 128 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=136120 $D=0
M2380 757 739 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=140750 $D=0
M2381 758 740 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=145380 $D=0
M2382 759 744 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=136120 $D=0
M2383 760 745 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=140750 $D=0
M2384 761 746 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=145380 $D=0
M2385 762 744 756 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=136120 $D=0
M2386 763 745 757 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=140750 $D=0
M2387 764 746 758 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=145380 $D=0
M2388 124 759 762 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=136120 $D=0
M2389 125 760 763 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=140750 $D=0
M2390 126 761 764 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=145380 $D=0
M2391 1062 727 7 7 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=135760 $D=0
M2392 1063 728 7 7 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=140390 $D=0
M2393 1064 729 7 7 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=145020 $D=0
M2394 765 124 1062 7 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=135760 $D=0
M2395 766 125 1063 7 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=140390 $D=0
M2396 767 126 1064 7 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=145020 $D=0
M2397 768 762 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=136120 $D=0
M2398 769 763 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=140750 $D=0
M2399 770 764 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=145380 $D=0
M2400 771 727 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=136120 $D=0
M2401 772 728 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=140750 $D=0
M2402 773 729 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=145380 $D=0
M2403 7 124 771 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=136120 $D=0
M2404 7 125 772 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=140750 $D=0
M2405 7 126 773 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=145380 $D=0
M2406 774 727 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=136120 $D=0
M2407 775 728 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=140750 $D=0
M2408 776 729 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=145380 $D=0
M2409 7 124 774 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=136120 $D=0
M2410 7 125 775 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=140750 $D=0
M2411 7 126 776 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=145380 $D=0
M2412 1065 727 7 7 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=135940 $D=0
M2413 1066 728 7 7 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=140570 $D=0
M2414 1067 729 7 7 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=145200 $D=0
M2415 780 124 1065 7 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=135940 $D=0
M2416 781 125 1066 7 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=140570 $D=0
M2417 782 126 1067 7 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=145200 $D=0
M2418 7 774 780 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=136120 $D=0
M2419 7 775 781 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=140750 $D=0
M2420 7 776 782 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=145380 $D=0
M2421 783 135 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=136120 $D=0
M2422 784 135 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=140750 $D=0
M2423 785 135 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=145380 $D=0
M2424 786 135 765 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=136120 $D=0
M2425 787 135 766 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=140750 $D=0
M2426 788 135 767 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=145380 $D=0
M2427 771 783 786 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=136120 $D=0
M2428 772 784 787 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=140750 $D=0
M2429 773 785 788 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=145380 $D=0
M2430 789 135 768 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=136120 $D=0
M2431 790 135 769 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=140750 $D=0
M2432 791 135 770 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=145380 $D=0
M2433 780 783 789 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=136120 $D=0
M2434 781 784 790 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=140750 $D=0
M2435 782 785 791 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=145380 $D=0
M2436 792 136 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=136120 $D=0
M2437 793 136 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=140750 $D=0
M2438 794 136 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=145380 $D=0
M2439 795 136 789 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=136120 $D=0
M2440 796 136 790 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=140750 $D=0
M2441 797 136 791 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=145380 $D=0
M2442 786 792 795 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=136120 $D=0
M2443 787 793 796 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=140750 $D=0
M2444 788 794 797 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=145380 $D=0
M2445 14 795 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=136120 $D=0
M2446 15 796 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=140750 $D=0
M2447 16 797 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=145380 $D=0
M2448 798 137 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=136120 $D=0
M2449 799 137 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=140750 $D=0
M2450 800 137 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=145380 $D=0
M2451 803 137 801 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=136120 $D=0
M2452 804 137 802 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=140750 $D=0
M2453 805 137 9 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=145380 $D=0
M2454 138 798 803 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=136120 $D=0
M2455 139 799 804 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=140750 $D=0
M2456 801 800 805 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=145380 $D=0
M2457 806 137 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=136120 $D=0
M2458 807 137 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=140750 $D=0
M2459 808 137 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=145380 $D=0
M2460 810 137 809 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=136120 $D=0
M2461 811 137 9 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=140750 $D=0
M2462 812 137 9 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=145380 $D=0
M2463 140 806 810 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=136120 $D=0
M2464 141 807 811 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=140750 $D=0
M2465 142 808 812 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=145380 $D=0
M2466 813 137 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=136120 $D=0
M2467 814 137 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=140750 $D=0
M2468 815 137 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=145380 $D=0
M2469 816 137 9 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=136120 $D=0
M2470 817 137 9 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=140750 $D=0
M2471 818 137 9 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=145380 $D=0
M2472 143 813 816 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=136120 $D=0
M2473 144 814 817 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=140750 $D=0
M2474 145 815 818 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=145380 $D=0
M2475 819 137 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=136120 $D=0
M2476 820 137 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=140750 $D=0
M2477 821 137 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=145380 $D=0
M2478 822 137 9 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=136120 $D=0
M2479 823 137 9 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=140750 $D=0
M2480 824 137 9 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=145380 $D=0
M2481 146 819 822 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=136120 $D=0
M2482 147 820 823 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=140750 $D=0
M2483 148 821 824 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=145380 $D=0
M2484 825 137 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=136120 $D=0
M2485 826 137 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=140750 $D=0
M2486 827 137 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=145380 $D=0
M2487 828 137 9 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=136120 $D=0
M2488 829 137 9 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=140750 $D=0
M2489 830 137 9 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=145380 $D=0
M2490 149 825 828 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=136120 $D=0
M2491 150 826 829 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=140750 $D=0
M2492 151 827 830 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=145380 $D=0
M2493 7 727 1047 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=136120 $D=0
M2494 7 728 1048 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=140750 $D=0
M2495 7 729 1049 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=145380 $D=0
M2496 139 1047 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=136120 $D=0
M2497 801 1048 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=140750 $D=0
M2498 802 1049 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=145380 $D=0
M2499 831 126 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=136120 $D=0
M2500 832 126 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=140750 $D=0
M2501 833 126 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=145380 $D=0
M2502 142 126 139 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=136120 $D=0
M2503 152 126 801 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=140750 $D=0
M2504 809 126 802 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=145380 $D=0
M2505 803 831 142 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=136120 $D=0
M2506 804 832 152 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=140750 $D=0
M2507 805 833 809 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=145380 $D=0
M2508 834 125 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=136120 $D=0
M2509 835 125 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=140750 $D=0
M2510 836 125 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=145380 $D=0
M2511 134 125 142 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=136120 $D=0
M2512 133 125 152 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=140750 $D=0
M2513 132 125 809 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=145380 $D=0
M2514 810 834 134 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=136120 $D=0
M2515 811 835 133 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=140750 $D=0
M2516 812 836 132 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=145380 $D=0
M2517 837 124 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=136120 $D=0
M2518 838 124 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=140750 $D=0
M2519 839 124 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=145380 $D=0
M2520 129 124 134 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=136120 $D=0
M2521 130 124 133 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=140750 $D=0
M2522 131 124 132 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=145380 $D=0
M2523 816 837 129 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=136120 $D=0
M2524 817 838 130 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=140750 $D=0
M2525 818 839 131 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=145380 $D=0
M2526 840 153 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=136120 $D=0
M2527 841 153 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=140750 $D=0
M2528 842 153 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=145380 $D=0
M2529 154 153 129 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=136120 $D=0
M2530 155 153 130 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=140750 $D=0
M2531 156 153 131 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=145380 $D=0
M2532 822 840 154 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=136120 $D=0
M2533 823 841 155 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=140750 $D=0
M2534 824 842 156 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=145380 $D=0
M2535 843 157 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=136120 $D=0
M2536 844 157 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=140750 $D=0
M2537 845 157 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=145380 $D=0
M2538 202 157 154 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=136120 $D=0
M2539 203 157 155 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=140750 $D=0
M2540 204 157 156 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=145380 $D=0
M2541 828 843 202 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=136120 $D=0
M2542 829 844 203 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=140750 $D=0
M2543 830 845 204 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=145380 $D=0
M2544 846 158 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=136120 $D=0
M2545 847 158 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=140750 $D=0
M2546 848 158 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=145380 $D=0
M2547 849 158 115 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=136120 $D=0
M2548 850 158 116 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=140750 $D=0
M2549 851 158 117 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=145380 $D=0
M2550 11 846 849 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=136120 $D=0
M2551 12 847 850 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=140750 $D=0
M2552 13 848 851 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=145380 $D=0
M2553 852 712 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=136120 $D=0
M2554 853 713 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=140750 $D=0
M2555 854 714 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=145380 $D=0
M2556 7 849 852 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=136120 $D=0
M2557 7 850 853 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=140750 $D=0
M2558 7 851 854 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=145380 $D=0
M2559 1068 712 7 7 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=135940 $D=0
M2560 1069 713 7 7 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=140570 $D=0
M2561 1070 714 7 7 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=145200 $D=0
M2562 858 849 1068 7 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=135940 $D=0
M2563 859 850 1069 7 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=140570 $D=0
M2564 860 851 1070 7 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=145200 $D=0
M2565 7 852 858 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=136120 $D=0
M2566 7 853 859 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=140750 $D=0
M2567 7 854 860 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=145380 $D=0
M2568 1050 159 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=136120 $D=0
M2569 1051 861 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=140750 $D=0
M2570 1052 862 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=145380 $D=0
M2571 7 858 1050 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=136120 $D=0
M2572 7 859 1051 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=140750 $D=0
M2573 7 860 1052 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=145380 $D=0
M2574 861 1050 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=136120 $D=0
M2575 862 1051 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=140750 $D=0
M2576 160 1052 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=145380 $D=0
M2577 1071 712 7 7 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=135760 $D=0
M2578 1072 713 7 7 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=140390 $D=0
M2579 1073 714 7 7 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=145020 $D=0
M2580 863 866 1071 7 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=135760 $D=0
M2581 864 867 1072 7 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=140390 $D=0
M2582 865 868 1073 7 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=145020 $D=0
M2583 866 849 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=136120 $D=0
M2584 867 850 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=140750 $D=0
M2585 868 851 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=145380 $D=0
M2586 869 863 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=136120 $D=0
M2587 870 864 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=140750 $D=0
M2588 871 865 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=145380 $D=0
M2589 7 159 869 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=136120 $D=0
M2590 7 861 870 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=140750 $D=0
M2591 7 862 871 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=145380 $D=0
M2592 874 161 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=136120 $D=0
M2593 875 872 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=140750 $D=0
M2594 876 873 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=145380 $D=0
M2595 872 869 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=136120 $D=0
M2596 873 870 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=140750 $D=0
M2597 162 871 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=145380 $D=0
M2598 7 874 872 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=136120 $D=0
M2599 7 875 873 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=140750 $D=0
M2600 7 876 162 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=145380 $D=0
M2601 879 877 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=136120 $D=0
M2602 880 878 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=140750 $D=0
M2603 881 9 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=145380 $D=0
M2604 7 885 882 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=136120 $D=0
M2605 7 886 883 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=140750 $D=0
M2606 7 887 884 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=145380 $D=0
M2607 888 119 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=136120 $D=0
M2608 889 120 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=140750 $D=0
M2609 890 121 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=145380 $D=0
M2610 885 119 877 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=136120 $D=0
M2611 886 120 878 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=140750 $D=0
M2612 887 121 9 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=145380 $D=0
M2613 879 888 885 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=136120 $D=0
M2614 880 889 886 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=140750 $D=0
M2615 881 890 887 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=145380 $D=0
M2616 891 882 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=136120 $D=0
M2617 892 883 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=140750 $D=0
M2618 893 884 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=145380 $D=0
M2619 163 882 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=136120 $D=0
M2620 877 883 9 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=140750 $D=0
M2621 878 884 9 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=145380 $D=0
M2622 119 891 163 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=136120 $D=0
M2623 120 892 877 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=140750 $D=0
M2624 121 893 878 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=145380 $D=0
M2625 894 163 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=136120 $D=0
M2626 895 877 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=140750 $D=0
M2627 896 878 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=145380 $D=0
M2628 897 882 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=136120 $D=0
M2629 898 883 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=140750 $D=0
M2630 899 884 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=145380 $D=0
M2631 205 882 894 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=136120 $D=0
M2632 206 883 895 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=140750 $D=0
M2633 207 884 896 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=145380 $D=0
M2634 7 897 205 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=136120 $D=0
M2635 9 898 206 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=140750 $D=0
M2636 9 899 207 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=145380 $D=0
M2637 900 164 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=136120 $D=0
M2638 901 164 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=140750 $D=0
M2639 902 164 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=145380 $D=0
M2640 903 164 205 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=136120 $D=0
M2641 904 164 206 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=140750 $D=0
M2642 905 164 207 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=145380 $D=0
M2643 14 900 903 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=136120 $D=0
M2644 15 901 904 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=140750 $D=0
M2645 16 902 905 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=145380 $D=0
M2646 906 165 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=136120 $D=0
M2647 907 165 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=140750 $D=0
M2648 908 165 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=145380 $D=0
M2649 909 165 903 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=136120 $D=0
M2650 910 165 904 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=140750 $D=0
M2651 911 165 905 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=145380 $D=0
M2652 9 906 909 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=136120 $D=0
M2653 9 907 910 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=140750 $D=0
M2654 9 908 911 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=145380 $D=0
M2655 912 114 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=136120 $D=0
M2656 913 114 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=140750 $D=0
M2657 914 114 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=145380 $D=0
M2658 7 912 915 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=136120 $D=0
M2659 7 913 916 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=140750 $D=0
M2660 7 914 917 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=145380 $D=0
M2661 918 114 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=136120 $D=0
M2662 919 114 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=140750 $D=0
M2663 920 114 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=145380 $D=0
M2664 921 915 909 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=136120 $D=0
M2665 922 916 910 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=140750 $D=0
M2666 923 917 911 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=145380 $D=0
M2667 7 921 1053 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=136120 $D=0
M2668 7 922 1054 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=140750 $D=0
M2669 7 923 1055 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=145380 $D=0
M2670 924 1053 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=136120 $D=0
M2671 925 1054 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=140750 $D=0
M2672 926 1055 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=145380 $D=0
M2673 921 912 924 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=136120 $D=0
M2674 922 913 925 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=140750 $D=0
M2675 923 914 926 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=145380 $D=0
M2676 927 918 924 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=136120 $D=0
M2677 928 919 925 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=140750 $D=0
M2678 929 920 926 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=145380 $D=0
M2679 7 933 930 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=136120 $D=0
M2680 7 934 931 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=140750 $D=0
M2681 7 935 932 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=145380 $D=0
M2682 933 114 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=136120 $D=0
M2683 934 114 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=140750 $D=0
M2684 935 114 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=145380 $D=0
M2685 1056 927 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=136120 $D=0
M2686 1057 928 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=140750 $D=0
M2687 1058 929 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=145380 $D=0
M2688 936 933 1056 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=136120 $D=0
M2689 937 934 1057 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=140750 $D=0
M2690 938 935 1058 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=145380 $D=0
M2691 7 936 119 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=136120 $D=0
M2692 7 937 120 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=140750 $D=0
M2693 7 938 121 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=145380 $D=0
M2694 1059 119 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=136120 $D=0
M2695 1060 120 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=140750 $D=0
M2696 1061 121 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=145380 $D=0
M2697 936 930 1059 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=136120 $D=0
M2698 937 931 1060 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=140750 $D=0
M2699 938 932 1061 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=145380 $D=0
.ENDS
***************************************
.SUBCKT ICV_25 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141
+ 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
** N=789 EP=159 IP=1514 FDC=1800
M0 176 1 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=125610 $D=1
M1 177 1 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=130240 $D=1
M2 178 176 2 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=125610 $D=1
M3 179 177 3 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=130240 $D=1
M4 8 1 178 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=125610 $D=1
M5 8 1 179 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=130240 $D=1
M6 180 176 2 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=125610 $D=1
M7 181 177 3 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=130240 $D=1
M8 2 1 180 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=125610 $D=1
M9 3 1 181 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=130240 $D=1
M10 182 176 2 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=125610 $D=1
M11 183 177 3 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=130240 $D=1
M12 2 1 182 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=125610 $D=1
M13 3 1 183 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=130240 $D=1
M14 186 184 182 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=125610 $D=1
M15 187 185 183 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=130240 $D=1
M16 184 4 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=125610 $D=1
M17 185 4 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=130240 $D=1
M18 188 184 180 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=125610 $D=1
M19 189 185 181 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=130240 $D=1
M20 178 4 188 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=125610 $D=1
M21 179 4 189 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=130240 $D=1
M22 190 5 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=125610 $D=1
M23 191 5 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=130240 $D=1
M24 192 190 188 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=125610 $D=1
M25 193 191 189 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=130240 $D=1
M26 186 5 192 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=125610 $D=1
M27 187 5 193 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=130240 $D=1
M28 194 7 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=125610 $D=1
M29 195 7 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=130240 $D=1
M30 196 194 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=125610 $D=1
M31 197 195 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=130240 $D=1
M32 9 7 196 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=125610 $D=1
M33 10 7 197 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=130240 $D=1
M34 198 194 11 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=125610 $D=1
M35 199 195 12 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=130240 $D=1
M36 200 7 198 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=125610 $D=1
M37 201 7 199 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=130240 $D=1
M38 204 194 202 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=125610 $D=1
M39 205 195 203 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=130240 $D=1
M40 192 7 204 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=125610 $D=1
M41 193 7 205 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=130240 $D=1
M42 208 206 204 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=125610 $D=1
M43 209 207 205 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=130240 $D=1
M44 206 13 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=125610 $D=1
M45 207 13 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=130240 $D=1
M46 210 206 198 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=125610 $D=1
M47 211 207 199 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=130240 $D=1
M48 196 13 210 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=125610 $D=1
M49 197 13 211 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=130240 $D=1
M50 212 14 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=125610 $D=1
M51 213 14 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=130240 $D=1
M52 214 212 210 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=125610 $D=1
M53 215 213 211 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=130240 $D=1
M54 208 14 214 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=125610 $D=1
M55 209 14 215 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=130240 $D=1
M56 8 15 216 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=125610 $D=1
M57 8 15 217 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=130240 $D=1
M58 218 16 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=125610 $D=1
M59 219 16 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=130240 $D=1
M60 220 15 214 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=125610 $D=1
M61 221 15 215 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=130240 $D=1
M62 8 220 688 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=125610 $D=1
M63 8 221 689 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=130240 $D=1
M64 222 688 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=125610 $D=1
M65 223 689 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=130240 $D=1
M66 220 216 222 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=125610 $D=1
M67 221 217 223 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=130240 $D=1
M68 222 16 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=125610 $D=1
M69 223 16 225 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=130240 $D=1
M70 228 17 222 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=125610 $D=1
M71 229 17 223 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=130240 $D=1
M72 226 17 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=125610 $D=1
M73 227 17 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=130240 $D=1
M74 8 18 230 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=125610 $D=1
M75 8 18 231 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=130240 $D=1
M76 232 19 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=125610 $D=1
M77 233 19 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=130240 $D=1
M78 234 18 214 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=125610 $D=1
M79 235 18 215 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=130240 $D=1
M80 8 234 690 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=125610 $D=1
M81 8 235 691 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=130240 $D=1
M82 236 690 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=125610 $D=1
M83 237 691 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=130240 $D=1
M84 234 230 236 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=125610 $D=1
M85 235 231 237 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=130240 $D=1
M86 236 19 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=125610 $D=1
M87 237 19 225 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=130240 $D=1
M88 228 20 236 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=125610 $D=1
M89 229 20 237 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=130240 $D=1
M90 238 20 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=125610 $D=1
M91 239 20 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=130240 $D=1
M92 8 21 240 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=125610 $D=1
M93 8 21 241 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=130240 $D=1
M94 242 22 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=125610 $D=1
M95 243 22 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=130240 $D=1
M96 244 21 214 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=125610 $D=1
M97 245 21 215 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=130240 $D=1
M98 8 244 692 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=125610 $D=1
M99 8 245 693 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=130240 $D=1
M100 246 692 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=125610 $D=1
M101 247 693 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=130240 $D=1
M102 244 240 246 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=125610 $D=1
M103 245 241 247 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=130240 $D=1
M104 246 22 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=125610 $D=1
M105 247 22 225 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=130240 $D=1
M106 228 23 246 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=125610 $D=1
M107 229 23 247 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=130240 $D=1
M108 248 23 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=125610 $D=1
M109 249 23 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=130240 $D=1
M110 8 24 250 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=125610 $D=1
M111 8 24 251 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=130240 $D=1
M112 252 25 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=125610 $D=1
M113 253 25 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=130240 $D=1
M114 254 24 214 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=125610 $D=1
M115 255 24 215 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=130240 $D=1
M116 8 254 694 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=125610 $D=1
M117 8 255 695 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=130240 $D=1
M118 256 694 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=125610 $D=1
M119 257 695 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=130240 $D=1
M120 254 250 256 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=125610 $D=1
M121 255 251 257 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=130240 $D=1
M122 256 25 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=125610 $D=1
M123 257 25 225 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=130240 $D=1
M124 228 26 256 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=125610 $D=1
M125 229 26 257 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=130240 $D=1
M126 258 26 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=125610 $D=1
M127 259 26 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=130240 $D=1
M128 8 27 260 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=125610 $D=1
M129 8 27 261 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=130240 $D=1
M130 262 28 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=125610 $D=1
M131 263 28 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=130240 $D=1
M132 264 27 214 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=125610 $D=1
M133 265 27 215 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=130240 $D=1
M134 8 264 696 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=125610 $D=1
M135 8 265 697 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=130240 $D=1
M136 266 696 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=125610 $D=1
M137 267 697 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=130240 $D=1
M138 264 260 266 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=125610 $D=1
M139 265 261 267 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=130240 $D=1
M140 266 28 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=125610 $D=1
M141 267 28 225 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=130240 $D=1
M142 228 29 266 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=125610 $D=1
M143 229 29 267 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=130240 $D=1
M144 268 29 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=125610 $D=1
M145 269 29 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=130240 $D=1
M146 8 30 270 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=125610 $D=1
M147 8 30 271 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=130240 $D=1
M148 272 31 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=125610 $D=1
M149 273 31 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=130240 $D=1
M150 274 30 214 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=125610 $D=1
M151 275 30 215 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=130240 $D=1
M152 8 274 698 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=125610 $D=1
M153 8 275 699 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=130240 $D=1
M154 276 698 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=125610 $D=1
M155 277 699 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=130240 $D=1
M156 274 270 276 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=125610 $D=1
M157 275 271 277 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=130240 $D=1
M158 276 31 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=125610 $D=1
M159 277 31 225 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=130240 $D=1
M160 228 32 276 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=125610 $D=1
M161 229 32 277 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=130240 $D=1
M162 278 32 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=125610 $D=1
M163 279 32 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=130240 $D=1
M164 8 33 280 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=125610 $D=1
M165 8 33 281 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=130240 $D=1
M166 282 34 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=125610 $D=1
M167 283 34 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=130240 $D=1
M168 284 33 214 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=125610 $D=1
M169 285 33 215 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=130240 $D=1
M170 8 284 700 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=125610 $D=1
M171 8 285 701 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=130240 $D=1
M172 286 700 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=125610 $D=1
M173 287 701 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=130240 $D=1
M174 284 280 286 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=125610 $D=1
M175 285 281 287 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=130240 $D=1
M176 286 34 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=125610 $D=1
M177 287 34 225 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=130240 $D=1
M178 228 35 286 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=125610 $D=1
M179 229 35 287 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=130240 $D=1
M180 288 35 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=125610 $D=1
M181 289 35 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=130240 $D=1
M182 8 36 290 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=125610 $D=1
M183 8 36 291 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=130240 $D=1
M184 292 37 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=125610 $D=1
M185 293 37 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=130240 $D=1
M186 294 36 214 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=125610 $D=1
M187 295 36 215 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=130240 $D=1
M188 8 294 702 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=125610 $D=1
M189 8 295 703 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=130240 $D=1
M190 296 702 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=125610 $D=1
M191 297 703 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=130240 $D=1
M192 294 290 296 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=125610 $D=1
M193 295 291 297 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=130240 $D=1
M194 296 37 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=125610 $D=1
M195 297 37 225 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=130240 $D=1
M196 228 38 296 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=125610 $D=1
M197 229 38 297 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=130240 $D=1
M198 298 38 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=125610 $D=1
M199 299 38 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=130240 $D=1
M200 8 39 300 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=125610 $D=1
M201 8 39 301 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=130240 $D=1
M202 302 40 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=125610 $D=1
M203 303 40 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=130240 $D=1
M204 304 39 214 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=125610 $D=1
M205 305 39 215 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=130240 $D=1
M206 8 304 704 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=125610 $D=1
M207 8 305 705 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=130240 $D=1
M208 306 704 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=125610 $D=1
M209 307 705 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=130240 $D=1
M210 304 300 306 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=125610 $D=1
M211 305 301 307 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=130240 $D=1
M212 306 40 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=125610 $D=1
M213 307 40 225 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=130240 $D=1
M214 228 41 306 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=125610 $D=1
M215 229 41 307 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=130240 $D=1
M216 308 41 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=125610 $D=1
M217 309 41 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=130240 $D=1
M218 8 42 310 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=125610 $D=1
M219 8 42 311 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=130240 $D=1
M220 312 43 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=125610 $D=1
M221 313 43 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=130240 $D=1
M222 314 42 214 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=125610 $D=1
M223 315 42 215 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=130240 $D=1
M224 8 314 706 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=125610 $D=1
M225 8 315 707 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=130240 $D=1
M226 316 706 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=125610 $D=1
M227 317 707 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=130240 $D=1
M228 314 310 316 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=125610 $D=1
M229 315 311 317 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=130240 $D=1
M230 316 43 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=125610 $D=1
M231 317 43 225 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=130240 $D=1
M232 228 44 316 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=125610 $D=1
M233 229 44 317 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=130240 $D=1
M234 318 44 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=125610 $D=1
M235 319 44 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=130240 $D=1
M236 8 45 320 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=125610 $D=1
M237 8 45 321 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=130240 $D=1
M238 322 46 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=125610 $D=1
M239 323 46 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=130240 $D=1
M240 324 45 214 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=125610 $D=1
M241 325 45 215 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=130240 $D=1
M242 8 324 708 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=125610 $D=1
M243 8 325 709 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=130240 $D=1
M244 326 708 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=125610 $D=1
M245 327 709 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=130240 $D=1
M246 324 320 326 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=125610 $D=1
M247 325 321 327 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=130240 $D=1
M248 326 46 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=125610 $D=1
M249 327 46 225 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=130240 $D=1
M250 228 47 326 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=125610 $D=1
M251 229 47 327 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=130240 $D=1
M252 328 47 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=125610 $D=1
M253 329 47 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=130240 $D=1
M254 8 48 330 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=125610 $D=1
M255 8 48 331 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=130240 $D=1
M256 332 49 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=125610 $D=1
M257 333 49 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=130240 $D=1
M258 334 48 214 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=125610 $D=1
M259 335 48 215 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=130240 $D=1
M260 8 334 710 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=125610 $D=1
M261 8 335 711 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=130240 $D=1
M262 336 710 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=125610 $D=1
M263 337 711 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=130240 $D=1
M264 334 330 336 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=125610 $D=1
M265 335 331 337 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=130240 $D=1
M266 336 49 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=125610 $D=1
M267 337 49 225 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=130240 $D=1
M268 228 50 336 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=125610 $D=1
M269 229 50 337 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=130240 $D=1
M270 338 50 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=125610 $D=1
M271 339 50 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=130240 $D=1
M272 8 51 340 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=125610 $D=1
M273 8 51 341 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=130240 $D=1
M274 342 52 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=125610 $D=1
M275 343 52 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=130240 $D=1
M276 344 51 214 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=125610 $D=1
M277 345 51 215 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=130240 $D=1
M278 8 344 712 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=125610 $D=1
M279 8 345 713 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=130240 $D=1
M280 346 712 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=125610 $D=1
M281 347 713 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=130240 $D=1
M282 344 340 346 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=125610 $D=1
M283 345 341 347 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=130240 $D=1
M284 346 52 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=125610 $D=1
M285 347 52 225 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=130240 $D=1
M286 228 53 346 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=125610 $D=1
M287 229 53 347 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=130240 $D=1
M288 348 53 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=125610 $D=1
M289 349 53 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=130240 $D=1
M290 8 54 350 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=125610 $D=1
M291 8 54 351 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=130240 $D=1
M292 352 55 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=125610 $D=1
M293 353 55 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=130240 $D=1
M294 354 54 214 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=125610 $D=1
M295 355 54 215 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=130240 $D=1
M296 8 354 714 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=125610 $D=1
M297 8 355 715 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=130240 $D=1
M298 356 714 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=125610 $D=1
M299 357 715 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=130240 $D=1
M300 354 350 356 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=125610 $D=1
M301 355 351 357 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=130240 $D=1
M302 356 55 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=125610 $D=1
M303 357 55 225 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=130240 $D=1
M304 228 56 356 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=125610 $D=1
M305 229 56 357 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=130240 $D=1
M306 358 56 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=125610 $D=1
M307 359 56 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=130240 $D=1
M308 8 57 360 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=125610 $D=1
M309 8 57 361 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=130240 $D=1
M310 362 58 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=125610 $D=1
M311 363 58 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=130240 $D=1
M312 364 57 214 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=125610 $D=1
M313 365 57 215 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=130240 $D=1
M314 8 364 716 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=125610 $D=1
M315 8 365 717 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=130240 $D=1
M316 366 716 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=125610 $D=1
M317 367 717 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=130240 $D=1
M318 364 360 366 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=125610 $D=1
M319 365 361 367 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=130240 $D=1
M320 366 58 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=125610 $D=1
M321 367 58 225 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=130240 $D=1
M322 228 59 366 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=125610 $D=1
M323 229 59 367 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=130240 $D=1
M324 368 59 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=125610 $D=1
M325 369 59 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=130240 $D=1
M326 8 60 370 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=125610 $D=1
M327 8 60 371 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=130240 $D=1
M328 372 61 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=125610 $D=1
M329 373 61 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=130240 $D=1
M330 374 60 214 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=125610 $D=1
M331 375 60 215 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=130240 $D=1
M332 8 374 718 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=125610 $D=1
M333 8 375 719 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=130240 $D=1
M334 376 718 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=125610 $D=1
M335 377 719 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=130240 $D=1
M336 374 370 376 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=125610 $D=1
M337 375 371 377 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=130240 $D=1
M338 376 61 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=125610 $D=1
M339 377 61 225 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=130240 $D=1
M340 228 62 376 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=125610 $D=1
M341 229 62 377 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=130240 $D=1
M342 378 62 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=125610 $D=1
M343 379 62 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=130240 $D=1
M344 8 63 380 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=125610 $D=1
M345 8 63 381 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=130240 $D=1
M346 382 64 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=125610 $D=1
M347 383 64 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=130240 $D=1
M348 384 63 214 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=125610 $D=1
M349 385 63 215 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=130240 $D=1
M350 8 384 720 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=125610 $D=1
M351 8 385 721 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=130240 $D=1
M352 386 720 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=125610 $D=1
M353 387 721 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=130240 $D=1
M354 384 380 386 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=125610 $D=1
M355 385 381 387 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=130240 $D=1
M356 386 64 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=125610 $D=1
M357 387 64 225 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=130240 $D=1
M358 228 65 386 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=125610 $D=1
M359 229 65 387 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=130240 $D=1
M360 388 65 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=125610 $D=1
M361 389 65 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=130240 $D=1
M362 8 66 390 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=125610 $D=1
M363 8 66 391 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=130240 $D=1
M364 392 67 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=125610 $D=1
M365 393 67 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=130240 $D=1
M366 394 66 214 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=125610 $D=1
M367 395 66 215 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=130240 $D=1
M368 8 394 722 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=125610 $D=1
M369 8 395 723 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=130240 $D=1
M370 396 722 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=125610 $D=1
M371 397 723 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=130240 $D=1
M372 394 390 396 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=125610 $D=1
M373 395 391 397 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=130240 $D=1
M374 396 67 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=125610 $D=1
M375 397 67 225 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=130240 $D=1
M376 228 68 396 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=125610 $D=1
M377 229 68 397 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=130240 $D=1
M378 398 68 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=125610 $D=1
M379 399 68 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=130240 $D=1
M380 8 69 400 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=125610 $D=1
M381 8 69 401 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=130240 $D=1
M382 402 70 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=125610 $D=1
M383 403 70 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=130240 $D=1
M384 404 69 214 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=125610 $D=1
M385 405 69 215 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=130240 $D=1
M386 8 404 724 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=125610 $D=1
M387 8 405 725 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=130240 $D=1
M388 406 724 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=125610 $D=1
M389 407 725 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=130240 $D=1
M390 404 400 406 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=125610 $D=1
M391 405 401 407 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=130240 $D=1
M392 406 70 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=125610 $D=1
M393 407 70 225 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=130240 $D=1
M394 228 71 406 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=125610 $D=1
M395 229 71 407 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=130240 $D=1
M396 408 71 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=125610 $D=1
M397 409 71 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=130240 $D=1
M398 8 72 410 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=125610 $D=1
M399 8 72 411 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=130240 $D=1
M400 412 73 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=125610 $D=1
M401 413 73 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=130240 $D=1
M402 414 72 214 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=125610 $D=1
M403 415 72 215 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=130240 $D=1
M404 8 414 726 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=125610 $D=1
M405 8 415 727 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=130240 $D=1
M406 416 726 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=125610 $D=1
M407 417 727 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=130240 $D=1
M408 414 410 416 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=125610 $D=1
M409 415 411 417 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=130240 $D=1
M410 416 73 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=125610 $D=1
M411 417 73 225 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=130240 $D=1
M412 228 74 416 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=125610 $D=1
M413 229 74 417 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=130240 $D=1
M414 418 74 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=125610 $D=1
M415 419 74 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=130240 $D=1
M416 8 75 420 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=125610 $D=1
M417 8 75 421 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=130240 $D=1
M418 422 76 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=125610 $D=1
M419 423 76 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=130240 $D=1
M420 424 75 214 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=125610 $D=1
M421 425 75 215 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=130240 $D=1
M422 8 424 728 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=125610 $D=1
M423 8 425 729 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=130240 $D=1
M424 426 728 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=125610 $D=1
M425 427 729 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=130240 $D=1
M426 424 420 426 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=125610 $D=1
M427 425 421 427 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=130240 $D=1
M428 426 76 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=125610 $D=1
M429 427 76 225 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=130240 $D=1
M430 228 77 426 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=125610 $D=1
M431 229 77 427 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=130240 $D=1
M432 428 77 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=125610 $D=1
M433 429 77 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=130240 $D=1
M434 8 78 430 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=125610 $D=1
M435 8 78 431 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=130240 $D=1
M436 432 79 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=125610 $D=1
M437 433 79 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=130240 $D=1
M438 434 78 214 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=125610 $D=1
M439 435 78 215 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=130240 $D=1
M440 8 434 730 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=125610 $D=1
M441 8 435 731 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=130240 $D=1
M442 436 730 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=125610 $D=1
M443 437 731 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=130240 $D=1
M444 434 430 436 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=125610 $D=1
M445 435 431 437 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=130240 $D=1
M446 436 79 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=125610 $D=1
M447 437 79 225 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=130240 $D=1
M448 228 80 436 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=125610 $D=1
M449 229 80 437 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=130240 $D=1
M450 438 80 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=125610 $D=1
M451 439 80 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=130240 $D=1
M452 8 81 440 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=125610 $D=1
M453 8 81 441 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=130240 $D=1
M454 442 82 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=125610 $D=1
M455 443 82 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=130240 $D=1
M456 444 81 214 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=125610 $D=1
M457 445 81 215 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=130240 $D=1
M458 8 444 732 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=125610 $D=1
M459 8 445 733 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=130240 $D=1
M460 446 732 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=125610 $D=1
M461 447 733 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=130240 $D=1
M462 444 440 446 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=125610 $D=1
M463 445 441 447 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=130240 $D=1
M464 446 82 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=125610 $D=1
M465 447 82 225 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=130240 $D=1
M466 228 83 446 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=125610 $D=1
M467 229 83 447 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=130240 $D=1
M468 448 83 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=125610 $D=1
M469 449 83 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=130240 $D=1
M470 8 84 450 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=125610 $D=1
M471 8 84 451 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=130240 $D=1
M472 452 85 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=125610 $D=1
M473 453 85 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=130240 $D=1
M474 454 84 214 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=125610 $D=1
M475 455 84 215 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=130240 $D=1
M476 8 454 734 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=125610 $D=1
M477 8 455 735 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=130240 $D=1
M478 456 734 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=125610 $D=1
M479 457 735 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=130240 $D=1
M480 454 450 456 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=125610 $D=1
M481 455 451 457 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=130240 $D=1
M482 456 85 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=125610 $D=1
M483 457 85 225 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=130240 $D=1
M484 228 86 456 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=125610 $D=1
M485 229 86 457 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=130240 $D=1
M486 458 86 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=125610 $D=1
M487 459 86 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=130240 $D=1
M488 8 87 460 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=125610 $D=1
M489 8 87 461 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=130240 $D=1
M490 462 88 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=125610 $D=1
M491 463 88 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=130240 $D=1
M492 464 87 214 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=125610 $D=1
M493 465 87 215 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=130240 $D=1
M494 8 464 736 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=125610 $D=1
M495 8 465 737 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=130240 $D=1
M496 466 736 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=125610 $D=1
M497 467 737 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=130240 $D=1
M498 464 460 466 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=125610 $D=1
M499 465 461 467 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=130240 $D=1
M500 466 88 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=125610 $D=1
M501 467 88 225 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=130240 $D=1
M502 228 89 466 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=125610 $D=1
M503 229 89 467 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=130240 $D=1
M504 468 89 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=125610 $D=1
M505 469 89 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=130240 $D=1
M506 8 90 470 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=125610 $D=1
M507 8 90 471 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=130240 $D=1
M508 472 91 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=125610 $D=1
M509 473 91 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=130240 $D=1
M510 474 90 214 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=125610 $D=1
M511 475 90 215 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=130240 $D=1
M512 8 474 738 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=125610 $D=1
M513 8 475 739 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=130240 $D=1
M514 476 738 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=125610 $D=1
M515 477 739 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=130240 $D=1
M516 474 470 476 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=125610 $D=1
M517 475 471 477 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=130240 $D=1
M518 476 91 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=125610 $D=1
M519 477 91 225 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=130240 $D=1
M520 228 92 476 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=125610 $D=1
M521 229 92 477 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=130240 $D=1
M522 478 92 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=125610 $D=1
M523 479 92 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=130240 $D=1
M524 8 93 480 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=125610 $D=1
M525 8 93 481 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=130240 $D=1
M526 482 94 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=125610 $D=1
M527 483 94 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=130240 $D=1
M528 484 93 214 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=125610 $D=1
M529 485 93 215 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=130240 $D=1
M530 8 484 740 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=125610 $D=1
M531 8 485 741 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=130240 $D=1
M532 486 740 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=125610 $D=1
M533 487 741 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=130240 $D=1
M534 484 480 486 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=125610 $D=1
M535 485 481 487 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=130240 $D=1
M536 486 94 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=125610 $D=1
M537 487 94 225 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=130240 $D=1
M538 228 95 486 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=125610 $D=1
M539 229 95 487 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=130240 $D=1
M540 488 95 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=125610 $D=1
M541 489 95 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=130240 $D=1
M542 8 96 490 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=125610 $D=1
M543 8 96 491 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=130240 $D=1
M544 492 97 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=125610 $D=1
M545 493 97 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=130240 $D=1
M546 494 96 214 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=125610 $D=1
M547 495 96 215 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=130240 $D=1
M548 8 494 742 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=125610 $D=1
M549 8 495 743 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=130240 $D=1
M550 496 742 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=125610 $D=1
M551 497 743 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=130240 $D=1
M552 494 490 496 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=125610 $D=1
M553 495 491 497 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=130240 $D=1
M554 496 97 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=125610 $D=1
M555 497 97 225 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=130240 $D=1
M556 228 98 496 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=125610 $D=1
M557 229 98 497 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=130240 $D=1
M558 498 98 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=125610 $D=1
M559 499 98 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=130240 $D=1
M560 8 99 500 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=125610 $D=1
M561 8 99 501 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=130240 $D=1
M562 502 100 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=125610 $D=1
M563 503 100 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=130240 $D=1
M564 504 99 214 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=125610 $D=1
M565 505 99 215 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=130240 $D=1
M566 8 504 744 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=125610 $D=1
M567 8 505 745 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=130240 $D=1
M568 506 744 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=125610 $D=1
M569 507 745 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=130240 $D=1
M570 504 500 506 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=125610 $D=1
M571 505 501 507 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=130240 $D=1
M572 506 100 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=125610 $D=1
M573 507 100 225 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=130240 $D=1
M574 228 101 506 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=125610 $D=1
M575 229 101 507 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=130240 $D=1
M576 508 101 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=125610 $D=1
M577 509 101 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=130240 $D=1
M578 8 102 510 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=125610 $D=1
M579 8 102 511 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=130240 $D=1
M580 512 103 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=125610 $D=1
M581 513 103 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=130240 $D=1
M582 514 102 214 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=125610 $D=1
M583 515 102 215 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=130240 $D=1
M584 8 514 746 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=125610 $D=1
M585 8 515 747 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=130240 $D=1
M586 516 746 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=125610 $D=1
M587 517 747 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=130240 $D=1
M588 514 510 516 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=125610 $D=1
M589 515 511 517 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=130240 $D=1
M590 516 103 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=125610 $D=1
M591 517 103 225 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=130240 $D=1
M592 228 104 516 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=125610 $D=1
M593 229 104 517 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=130240 $D=1
M594 518 104 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=125610 $D=1
M595 519 104 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=130240 $D=1
M596 8 105 520 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=125610 $D=1
M597 8 105 521 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=130240 $D=1
M598 522 106 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=125610 $D=1
M599 523 106 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=130240 $D=1
M600 524 105 214 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=125610 $D=1
M601 525 105 215 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=130240 $D=1
M602 8 524 748 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=125610 $D=1
M603 8 525 749 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=130240 $D=1
M604 526 748 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=125610 $D=1
M605 527 749 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=130240 $D=1
M606 524 520 526 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=125610 $D=1
M607 525 521 527 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=130240 $D=1
M608 526 106 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=125610 $D=1
M609 527 106 225 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=130240 $D=1
M610 228 107 526 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=125610 $D=1
M611 229 107 527 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=130240 $D=1
M612 528 107 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=125610 $D=1
M613 529 107 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=130240 $D=1
M614 8 108 530 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=125610 $D=1
M615 8 108 531 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=130240 $D=1
M616 532 109 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=125610 $D=1
M617 533 109 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=130240 $D=1
M618 8 109 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=125610 $D=1
M619 8 109 225 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=130240 $D=1
M620 228 108 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=125610 $D=1
M621 229 108 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=130240 $D=1
M622 8 536 534 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=125610 $D=1
M623 8 537 535 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=130240 $D=1
M624 536 110 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=125610 $D=1
M625 537 110 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=130240 $D=1
M626 750 224 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=125610 $D=1
M627 751 225 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=130240 $D=1
M628 538 534 750 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=125610 $D=1
M629 539 535 751 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=130240 $D=1
M630 8 538 540 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=125610 $D=1
M631 8 539 541 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=130240 $D=1
M632 752 540 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=125610 $D=1
M633 753 541 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=130240 $D=1
M634 538 536 752 8 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=125610 $D=1
M635 539 537 753 8 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=130240 $D=1
M636 8 544 542 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=125610 $D=1
M637 8 545 543 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=130240 $D=1
M638 544 110 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=125610 $D=1
M639 545 110 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=130240 $D=1
M640 754 228 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=125610 $D=1
M641 755 229 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=130240 $D=1
M642 546 542 754 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=125610 $D=1
M643 547 543 755 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=130240 $D=1
M644 8 546 111 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=125610 $D=1
M645 8 547 112 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=130240 $D=1
M646 756 111 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=125610 $D=1
M647 757 112 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=130240 $D=1
M648 546 544 756 8 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=125610 $D=1
M649 547 545 757 8 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=130240 $D=1
M650 548 113 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=125610 $D=1
M651 549 113 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=130240 $D=1
M652 550 548 540 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=125610 $D=1
M653 551 549 541 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=130240 $D=1
M654 114 113 550 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=125610 $D=1
M655 115 113 551 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=130240 $D=1
M656 552 116 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=125610 $D=1
M657 553 116 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=130240 $D=1
M658 554 552 111 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=125610 $D=1
M659 555 553 112 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=130240 $D=1
M660 758 116 554 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=125610 $D=1
M661 759 116 555 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=130240 $D=1
M662 8 111 758 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=125610 $D=1
M663 8 112 759 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=130240 $D=1
M664 556 117 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=125610 $D=1
M665 557 117 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=130240 $D=1
M666 118 556 554 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=125610 $D=1
M667 119 557 555 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=130240 $D=1
M668 9 117 118 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=125610 $D=1
M669 10 117 119 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=130240 $D=1
M670 559 558 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=125610 $D=1
M671 560 120 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=130240 $D=1
M672 8 563 561 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=125610 $D=1
M673 8 564 562 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=130240 $D=1
M674 565 550 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=125610 $D=1
M675 566 551 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=130240 $D=1
M676 563 565 558 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=125610 $D=1
M677 564 566 120 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=130240 $D=1
M678 559 550 563 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=125610 $D=1
M679 560 551 564 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=130240 $D=1
M680 567 561 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=125610 $D=1
M681 568 562 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=130240 $D=1
M682 121 567 118 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=125610 $D=1
M683 558 568 119 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=130240 $D=1
M684 550 561 121 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=125610 $D=1
M685 551 562 558 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=130240 $D=1
M686 569 121 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=125610 $D=1
M687 570 558 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=130240 $D=1
M688 571 561 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=125610 $D=1
M689 572 562 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=130240 $D=1
M690 573 571 569 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=125610 $D=1
M691 574 572 570 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=130240 $D=1
M692 118 561 573 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=125610 $D=1
M693 119 562 574 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=130240 $D=1
M694 575 550 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=125610 $D=1
M695 576 551 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=130240 $D=1
M696 8 118 575 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=125610 $D=1
M697 8 119 576 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=130240 $D=1
M698 577 573 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=125610 $D=1
M699 578 574 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=130240 $D=1
M700 778 550 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=125610 $D=1
M701 779 551 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=130240 $D=1
M702 579 118 778 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=125610 $D=1
M703 580 119 779 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=130240 $D=1
M704 780 550 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=125610 $D=1
M705 781 551 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=130240 $D=1
M706 581 118 780 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=125610 $D=1
M707 582 119 781 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=130240 $D=1
M708 585 550 583 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=125610 $D=1
M709 586 551 584 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=130240 $D=1
M710 583 118 585 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=125610 $D=1
M711 584 119 586 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=130240 $D=1
M712 8 581 583 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=125610 $D=1
M713 8 582 584 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=130240 $D=1
M714 587 127 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=125610 $D=1
M715 588 127 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=130240 $D=1
M716 589 587 575 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=125610 $D=1
M717 590 588 576 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=130240 $D=1
M718 579 127 589 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=125610 $D=1
M719 580 127 590 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=130240 $D=1
M720 591 587 577 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=125610 $D=1
M721 592 588 578 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=130240 $D=1
M722 585 127 591 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=125610 $D=1
M723 586 127 592 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=130240 $D=1
M724 593 128 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=125610 $D=1
M725 594 128 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=130240 $D=1
M726 595 593 591 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=125610 $D=1
M727 596 594 592 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=130240 $D=1
M728 589 128 595 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=125610 $D=1
M729 590 128 596 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=130240 $D=1
M730 11 595 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=125610 $D=1
M731 12 596 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=130240 $D=1
M732 597 130 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=125610 $D=1
M733 598 130 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=130240 $D=1
M734 599 597 131 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=125610 $D=1
M735 600 598 132 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=130240 $D=1
M736 133 130 599 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=125610 $D=1
M737 134 130 600 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=130240 $D=1
M738 601 130 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=125610 $D=1
M739 602 130 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=130240 $D=1
M740 603 601 135 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=125610 $D=1
M741 604 602 136 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=130240 $D=1
M742 137 130 603 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=125610 $D=1
M743 138 130 604 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=130240 $D=1
M744 605 130 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=125610 $D=1
M745 606 130 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=130240 $D=1
M746 607 605 124 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=125610 $D=1
M747 608 606 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=130240 $D=1
M748 129 130 607 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=125610 $D=1
M749 139 130 608 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=130240 $D=1
M750 609 130 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=125610 $D=1
M751 610 130 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=130240 $D=1
M752 611 609 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=125610 $D=1
M753 612 610 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=130240 $D=1
M754 140 130 611 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=125610 $D=1
M755 141 130 612 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=130240 $D=1
M756 613 130 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=125610 $D=1
M757 614 130 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=130240 $D=1
M758 615 613 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=125610 $D=1
M759 616 614 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=130240 $D=1
M760 142 130 615 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=125610 $D=1
M761 143 130 616 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=130240 $D=1
M762 8 550 760 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=125610 $D=1
M763 8 551 761 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=130240 $D=1
M764 134 760 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=125610 $D=1
M765 131 761 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=130240 $D=1
M766 617 144 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=125610 $D=1
M767 618 144 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=130240 $D=1
M768 145 617 134 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=125610 $D=1
M769 146 618 131 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=130240 $D=1
M770 599 144 145 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=125610 $D=1
M771 600 144 146 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=130240 $D=1
M772 619 147 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=125610 $D=1
M773 620 147 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=130240 $D=1
M774 148 619 145 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=125610 $D=1
M775 126 620 146 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=130240 $D=1
M776 603 147 148 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=125610 $D=1
M777 604 147 126 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=130240 $D=1
M778 621 149 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=125610 $D=1
M779 622 149 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=130240 $D=1
M780 122 621 148 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=125610 $D=1
M781 123 622 126 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=130240 $D=1
M782 607 149 122 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=125610 $D=1
M783 608 149 123 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=130240 $D=1
M784 623 119 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=125610 $D=1
M785 624 119 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=130240 $D=1
M786 150 623 122 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=125610 $D=1
M787 151 624 123 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=130240 $D=1
M788 611 119 150 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=125610 $D=1
M789 612 119 151 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=130240 $D=1
M790 625 118 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=125610 $D=1
M791 626 118 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=130240 $D=1
M792 200 625 150 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=125610 $D=1
M793 201 626 151 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=130240 $D=1
M794 615 118 200 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=125610 $D=1
M795 616 118 201 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=130240 $D=1
M796 627 152 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=125610 $D=1
M797 628 152 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=130240 $D=1
M798 629 627 111 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=125610 $D=1
M799 630 628 112 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=130240 $D=1
M800 9 152 629 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=125610 $D=1
M801 10 152 630 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=130240 $D=1
M802 782 540 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=125610 $D=1
M803 783 541 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=130240 $D=1
M804 631 629 782 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=125610 $D=1
M805 632 630 783 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=130240 $D=1
M806 635 540 633 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=125610 $D=1
M807 636 541 634 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=130240 $D=1
M808 633 629 635 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=125610 $D=1
M809 634 630 636 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=130240 $D=1
M810 8 631 633 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=125610 $D=1
M811 8 632 634 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=130240 $D=1
M812 784 153 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=125610 $D=1
M813 785 637 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=130240 $D=1
M814 762 635 784 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=125610 $D=1
M815 763 636 785 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=130240 $D=1
M816 637 762 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=125610 $D=1
M817 154 763 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=130240 $D=1
M818 638 540 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=125610 $D=1
M819 639 541 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=130240 $D=1
M820 8 640 638 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=125610 $D=1
M821 8 641 639 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=130240 $D=1
M822 640 629 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=125610 $D=1
M823 641 630 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=130240 $D=1
M824 786 638 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=125610 $D=1
M825 787 639 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=130240 $D=1
M826 642 153 786 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=125610 $D=1
M827 643 637 787 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=130240 $D=1
M828 645 155 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=125610 $D=1
M829 646 644 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=130240 $D=1
M830 788 642 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=125610 $D=1
M831 789 643 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=130240 $D=1
M832 644 645 788 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=125610 $D=1
M833 156 646 789 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=130240 $D=1
M834 648 647 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=125610 $D=1
M835 649 157 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=130240 $D=1
M836 8 652 650 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=125610 $D=1
M837 8 653 651 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=130240 $D=1
M838 654 114 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=125610 $D=1
M839 655 115 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=130240 $D=1
M840 652 654 647 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=125610 $D=1
M841 653 655 157 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=130240 $D=1
M842 648 114 652 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=125610 $D=1
M843 649 115 653 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=130240 $D=1
M844 656 650 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=125610 $D=1
M845 657 651 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=130240 $D=1
M846 158 656 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=125610 $D=1
M847 647 657 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=130240 $D=1
M848 114 650 158 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=125610 $D=1
M849 115 651 647 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=130240 $D=1
M850 658 158 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=125610 $D=1
M851 659 647 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=130240 $D=1
M852 660 650 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=125610 $D=1
M853 661 651 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=130240 $D=1
M854 202 660 658 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=125610 $D=1
M855 203 661 659 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=130240 $D=1
M856 8 650 202 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=125610 $D=1
M857 8 651 203 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=130240 $D=1
M858 662 159 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=125610 $D=1
M859 663 159 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=130240 $D=1
M860 664 662 202 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=125610 $D=1
M861 665 663 203 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=130240 $D=1
M862 11 159 664 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=125610 $D=1
M863 12 159 665 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=130240 $D=1
M864 666 160 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=125610 $D=1
M865 667 160 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=130240 $D=1
M866 668 666 664 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=125610 $D=1
M867 669 667 665 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=130240 $D=1
M868 8 160 668 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=125610 $D=1
M869 8 160 669 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=130240 $D=1
M870 670 110 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=125610 $D=1
M871 671 110 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=130240 $D=1
M872 8 670 672 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=125610 $D=1
M873 8 671 673 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=130240 $D=1
M874 674 110 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=125610 $D=1
M875 675 110 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=130240 $D=1
M876 676 670 668 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=125610 $D=1
M877 677 671 669 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=130240 $D=1
M878 8 676 764 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=125610 $D=1
M879 8 677 765 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=130240 $D=1
M880 678 764 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=125610 $D=1
M881 679 765 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=130240 $D=1
M882 676 672 678 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=125610 $D=1
M883 677 673 679 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=130240 $D=1
M884 680 110 678 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=125610 $D=1
M885 681 110 679 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=130240 $D=1
M886 8 684 682 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=125610 $D=1
M887 8 685 683 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=130240 $D=1
M888 684 110 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=125610 $D=1
M889 685 110 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=130240 $D=1
M890 766 680 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=125610 $D=1
M891 767 681 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=130240 $D=1
M892 686 682 766 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=125610 $D=1
M893 687 683 767 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=130240 $D=1
M894 8 686 114 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=125610 $D=1
M895 8 687 115 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=130240 $D=1
M896 768 114 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=125610 $D=1
M897 769 115 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=130240 $D=1
M898 686 684 768 8 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=125610 $D=1
M899 687 685 769 8 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=130240 $D=1
M900 176 1 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=126860 $D=0
M901 177 1 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=131490 $D=0
M902 178 1 2 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=126860 $D=0
M903 179 1 3 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=131490 $D=0
M904 8 176 178 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=126860 $D=0
M905 8 177 179 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=131490 $D=0
M906 180 1 2 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=126860 $D=0
M907 181 1 3 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=131490 $D=0
M908 2 176 180 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=126860 $D=0
M909 3 177 181 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=131490 $D=0
M910 182 1 2 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=126860 $D=0
M911 183 1 3 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=131490 $D=0
M912 2 176 182 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=126860 $D=0
M913 3 177 183 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=131490 $D=0
M914 186 4 182 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=126860 $D=0
M915 187 4 183 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=131490 $D=0
M916 184 4 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=126860 $D=0
M917 185 4 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=131490 $D=0
M918 188 4 180 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=126860 $D=0
M919 189 4 181 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=131490 $D=0
M920 178 184 188 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=126860 $D=0
M921 179 185 189 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=131490 $D=0
M922 190 5 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=126860 $D=0
M923 191 5 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=131490 $D=0
M924 192 5 188 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=126860 $D=0
M925 193 5 189 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=131490 $D=0
M926 186 190 192 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=126860 $D=0
M927 187 191 193 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=131490 $D=0
M928 194 7 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=126860 $D=0
M929 195 7 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=131490 $D=0
M930 196 7 8 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=126860 $D=0
M931 197 7 8 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=131490 $D=0
M932 9 194 196 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=126860 $D=0
M933 10 195 197 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=131490 $D=0
M934 198 7 11 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=126860 $D=0
M935 199 7 12 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=131490 $D=0
M936 200 194 198 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=126860 $D=0
M937 201 195 199 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=131490 $D=0
M938 204 7 202 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=126860 $D=0
M939 205 7 203 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=131490 $D=0
M940 192 194 204 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=126860 $D=0
M941 193 195 205 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=131490 $D=0
M942 208 13 204 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=126860 $D=0
M943 209 13 205 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=131490 $D=0
M944 206 13 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=126860 $D=0
M945 207 13 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=131490 $D=0
M946 210 13 198 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=126860 $D=0
M947 211 13 199 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=131490 $D=0
M948 196 206 210 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=126860 $D=0
M949 197 207 211 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=131490 $D=0
M950 212 14 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=126860 $D=0
M951 213 14 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=131490 $D=0
M952 214 14 210 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=126860 $D=0
M953 215 14 211 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=131490 $D=0
M954 208 212 214 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=126860 $D=0
M955 209 213 215 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=131490 $D=0
M956 6 15 216 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=126860 $D=0
M957 6 15 217 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=131490 $D=0
M958 218 16 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=126860 $D=0
M959 219 16 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=131490 $D=0
M960 220 216 214 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=126860 $D=0
M961 221 217 215 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=131490 $D=0
M962 6 220 688 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=126860 $D=0
M963 6 221 689 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=131490 $D=0
M964 222 688 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=126860 $D=0
M965 223 689 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=131490 $D=0
M966 220 15 222 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=126860 $D=0
M967 221 15 223 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=131490 $D=0
M968 222 218 224 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=126860 $D=0
M969 223 219 225 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=131490 $D=0
M970 228 226 222 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=126860 $D=0
M971 229 227 223 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=131490 $D=0
M972 226 17 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=126860 $D=0
M973 227 17 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=131490 $D=0
M974 6 18 230 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=126860 $D=0
M975 6 18 231 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=131490 $D=0
M976 232 19 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=126860 $D=0
M977 233 19 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=131490 $D=0
M978 234 230 214 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=126860 $D=0
M979 235 231 215 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=131490 $D=0
M980 6 234 690 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=126860 $D=0
M981 6 235 691 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=131490 $D=0
M982 236 690 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=126860 $D=0
M983 237 691 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=131490 $D=0
M984 234 18 236 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=126860 $D=0
M985 235 18 237 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=131490 $D=0
M986 236 232 224 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=126860 $D=0
M987 237 233 225 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=131490 $D=0
M988 228 238 236 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=126860 $D=0
M989 229 239 237 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=131490 $D=0
M990 238 20 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=126860 $D=0
M991 239 20 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=131490 $D=0
M992 6 21 240 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=126860 $D=0
M993 6 21 241 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=131490 $D=0
M994 242 22 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=126860 $D=0
M995 243 22 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=131490 $D=0
M996 244 240 214 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=126860 $D=0
M997 245 241 215 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=131490 $D=0
M998 6 244 692 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=126860 $D=0
M999 6 245 693 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=131490 $D=0
M1000 246 692 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=126860 $D=0
M1001 247 693 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=131490 $D=0
M1002 244 21 246 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=126860 $D=0
M1003 245 21 247 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=131490 $D=0
M1004 246 242 224 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=126860 $D=0
M1005 247 243 225 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=131490 $D=0
M1006 228 248 246 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=126860 $D=0
M1007 229 249 247 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=131490 $D=0
M1008 248 23 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=126860 $D=0
M1009 249 23 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=131490 $D=0
M1010 6 24 250 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=126860 $D=0
M1011 6 24 251 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=131490 $D=0
M1012 252 25 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=126860 $D=0
M1013 253 25 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=131490 $D=0
M1014 254 250 214 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=126860 $D=0
M1015 255 251 215 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=131490 $D=0
M1016 6 254 694 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=126860 $D=0
M1017 6 255 695 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=131490 $D=0
M1018 256 694 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=126860 $D=0
M1019 257 695 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=131490 $D=0
M1020 254 24 256 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=126860 $D=0
M1021 255 24 257 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=131490 $D=0
M1022 256 252 224 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=126860 $D=0
M1023 257 253 225 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=131490 $D=0
M1024 228 258 256 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=126860 $D=0
M1025 229 259 257 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=131490 $D=0
M1026 258 26 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=126860 $D=0
M1027 259 26 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=131490 $D=0
M1028 6 27 260 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=126860 $D=0
M1029 6 27 261 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=131490 $D=0
M1030 262 28 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=126860 $D=0
M1031 263 28 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=131490 $D=0
M1032 264 260 214 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=126860 $D=0
M1033 265 261 215 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=131490 $D=0
M1034 6 264 696 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=126860 $D=0
M1035 6 265 697 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=131490 $D=0
M1036 266 696 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=126860 $D=0
M1037 267 697 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=131490 $D=0
M1038 264 27 266 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=126860 $D=0
M1039 265 27 267 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=131490 $D=0
M1040 266 262 224 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=126860 $D=0
M1041 267 263 225 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=131490 $D=0
M1042 228 268 266 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=126860 $D=0
M1043 229 269 267 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=131490 $D=0
M1044 268 29 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=126860 $D=0
M1045 269 29 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=131490 $D=0
M1046 6 30 270 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=126860 $D=0
M1047 6 30 271 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=131490 $D=0
M1048 272 31 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=126860 $D=0
M1049 273 31 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=131490 $D=0
M1050 274 270 214 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=126860 $D=0
M1051 275 271 215 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=131490 $D=0
M1052 6 274 698 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=126860 $D=0
M1053 6 275 699 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=131490 $D=0
M1054 276 698 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=126860 $D=0
M1055 277 699 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=131490 $D=0
M1056 274 30 276 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=126860 $D=0
M1057 275 30 277 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=131490 $D=0
M1058 276 272 224 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=126860 $D=0
M1059 277 273 225 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=131490 $D=0
M1060 228 278 276 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=126860 $D=0
M1061 229 279 277 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=131490 $D=0
M1062 278 32 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=126860 $D=0
M1063 279 32 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=131490 $D=0
M1064 6 33 280 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=126860 $D=0
M1065 6 33 281 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=131490 $D=0
M1066 282 34 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=126860 $D=0
M1067 283 34 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=131490 $D=0
M1068 284 280 214 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=126860 $D=0
M1069 285 281 215 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=131490 $D=0
M1070 6 284 700 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=126860 $D=0
M1071 6 285 701 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=131490 $D=0
M1072 286 700 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=126860 $D=0
M1073 287 701 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=131490 $D=0
M1074 284 33 286 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=126860 $D=0
M1075 285 33 287 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=131490 $D=0
M1076 286 282 224 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=126860 $D=0
M1077 287 283 225 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=131490 $D=0
M1078 228 288 286 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=126860 $D=0
M1079 229 289 287 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=131490 $D=0
M1080 288 35 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=126860 $D=0
M1081 289 35 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=131490 $D=0
M1082 6 36 290 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=126860 $D=0
M1083 6 36 291 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=131490 $D=0
M1084 292 37 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=126860 $D=0
M1085 293 37 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=131490 $D=0
M1086 294 290 214 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=126860 $D=0
M1087 295 291 215 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=131490 $D=0
M1088 6 294 702 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=126860 $D=0
M1089 6 295 703 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=131490 $D=0
M1090 296 702 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=126860 $D=0
M1091 297 703 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=131490 $D=0
M1092 294 36 296 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=126860 $D=0
M1093 295 36 297 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=131490 $D=0
M1094 296 292 224 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=126860 $D=0
M1095 297 293 225 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=131490 $D=0
M1096 228 298 296 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=126860 $D=0
M1097 229 299 297 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=131490 $D=0
M1098 298 38 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=126860 $D=0
M1099 299 38 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=131490 $D=0
M1100 6 39 300 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=126860 $D=0
M1101 6 39 301 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=131490 $D=0
M1102 302 40 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=126860 $D=0
M1103 303 40 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=131490 $D=0
M1104 304 300 214 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=126860 $D=0
M1105 305 301 215 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=131490 $D=0
M1106 6 304 704 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=126860 $D=0
M1107 6 305 705 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=131490 $D=0
M1108 306 704 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=126860 $D=0
M1109 307 705 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=131490 $D=0
M1110 304 39 306 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=126860 $D=0
M1111 305 39 307 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=131490 $D=0
M1112 306 302 224 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=126860 $D=0
M1113 307 303 225 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=131490 $D=0
M1114 228 308 306 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=126860 $D=0
M1115 229 309 307 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=131490 $D=0
M1116 308 41 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=126860 $D=0
M1117 309 41 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=131490 $D=0
M1118 6 42 310 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=126860 $D=0
M1119 6 42 311 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=131490 $D=0
M1120 312 43 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=126860 $D=0
M1121 313 43 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=131490 $D=0
M1122 314 310 214 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=126860 $D=0
M1123 315 311 215 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=131490 $D=0
M1124 6 314 706 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=126860 $D=0
M1125 6 315 707 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=131490 $D=0
M1126 316 706 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=126860 $D=0
M1127 317 707 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=131490 $D=0
M1128 314 42 316 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=126860 $D=0
M1129 315 42 317 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=131490 $D=0
M1130 316 312 224 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=126860 $D=0
M1131 317 313 225 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=131490 $D=0
M1132 228 318 316 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=126860 $D=0
M1133 229 319 317 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=131490 $D=0
M1134 318 44 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=126860 $D=0
M1135 319 44 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=131490 $D=0
M1136 6 45 320 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=126860 $D=0
M1137 6 45 321 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=131490 $D=0
M1138 322 46 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=126860 $D=0
M1139 323 46 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=131490 $D=0
M1140 324 320 214 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=126860 $D=0
M1141 325 321 215 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=131490 $D=0
M1142 6 324 708 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=126860 $D=0
M1143 6 325 709 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=131490 $D=0
M1144 326 708 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=126860 $D=0
M1145 327 709 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=131490 $D=0
M1146 324 45 326 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=126860 $D=0
M1147 325 45 327 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=131490 $D=0
M1148 326 322 224 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=126860 $D=0
M1149 327 323 225 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=131490 $D=0
M1150 228 328 326 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=126860 $D=0
M1151 229 329 327 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=131490 $D=0
M1152 328 47 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=126860 $D=0
M1153 329 47 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=131490 $D=0
M1154 6 48 330 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=126860 $D=0
M1155 6 48 331 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=131490 $D=0
M1156 332 49 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=126860 $D=0
M1157 333 49 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=131490 $D=0
M1158 334 330 214 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=126860 $D=0
M1159 335 331 215 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=131490 $D=0
M1160 6 334 710 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=126860 $D=0
M1161 6 335 711 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=131490 $D=0
M1162 336 710 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=126860 $D=0
M1163 337 711 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=131490 $D=0
M1164 334 48 336 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=126860 $D=0
M1165 335 48 337 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=131490 $D=0
M1166 336 332 224 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=126860 $D=0
M1167 337 333 225 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=131490 $D=0
M1168 228 338 336 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=126860 $D=0
M1169 229 339 337 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=131490 $D=0
M1170 338 50 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=126860 $D=0
M1171 339 50 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=131490 $D=0
M1172 6 51 340 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=126860 $D=0
M1173 6 51 341 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=131490 $D=0
M1174 342 52 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=126860 $D=0
M1175 343 52 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=131490 $D=0
M1176 344 340 214 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=126860 $D=0
M1177 345 341 215 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=131490 $D=0
M1178 6 344 712 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=126860 $D=0
M1179 6 345 713 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=131490 $D=0
M1180 346 712 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=126860 $D=0
M1181 347 713 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=131490 $D=0
M1182 344 51 346 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=126860 $D=0
M1183 345 51 347 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=131490 $D=0
M1184 346 342 224 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=126860 $D=0
M1185 347 343 225 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=131490 $D=0
M1186 228 348 346 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=126860 $D=0
M1187 229 349 347 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=131490 $D=0
M1188 348 53 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=126860 $D=0
M1189 349 53 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=131490 $D=0
M1190 6 54 350 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=126860 $D=0
M1191 6 54 351 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=131490 $D=0
M1192 352 55 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=126860 $D=0
M1193 353 55 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=131490 $D=0
M1194 354 350 214 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=126860 $D=0
M1195 355 351 215 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=131490 $D=0
M1196 6 354 714 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=126860 $D=0
M1197 6 355 715 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=131490 $D=0
M1198 356 714 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=126860 $D=0
M1199 357 715 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=131490 $D=0
M1200 354 54 356 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=126860 $D=0
M1201 355 54 357 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=131490 $D=0
M1202 356 352 224 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=126860 $D=0
M1203 357 353 225 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=131490 $D=0
M1204 228 358 356 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=126860 $D=0
M1205 229 359 357 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=131490 $D=0
M1206 358 56 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=126860 $D=0
M1207 359 56 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=131490 $D=0
M1208 6 57 360 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=126860 $D=0
M1209 6 57 361 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=131490 $D=0
M1210 362 58 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=126860 $D=0
M1211 363 58 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=131490 $D=0
M1212 364 360 214 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=126860 $D=0
M1213 365 361 215 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=131490 $D=0
M1214 6 364 716 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=126860 $D=0
M1215 6 365 717 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=131490 $D=0
M1216 366 716 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=126860 $D=0
M1217 367 717 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=131490 $D=0
M1218 364 57 366 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=126860 $D=0
M1219 365 57 367 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=131490 $D=0
M1220 366 362 224 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=126860 $D=0
M1221 367 363 225 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=131490 $D=0
M1222 228 368 366 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=126860 $D=0
M1223 229 369 367 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=131490 $D=0
M1224 368 59 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=126860 $D=0
M1225 369 59 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=131490 $D=0
M1226 6 60 370 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=126860 $D=0
M1227 6 60 371 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=131490 $D=0
M1228 372 61 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=126860 $D=0
M1229 373 61 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=131490 $D=0
M1230 374 370 214 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=126860 $D=0
M1231 375 371 215 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=131490 $D=0
M1232 6 374 718 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=126860 $D=0
M1233 6 375 719 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=131490 $D=0
M1234 376 718 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=126860 $D=0
M1235 377 719 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=131490 $D=0
M1236 374 60 376 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=126860 $D=0
M1237 375 60 377 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=131490 $D=0
M1238 376 372 224 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=126860 $D=0
M1239 377 373 225 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=131490 $D=0
M1240 228 378 376 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=126860 $D=0
M1241 229 379 377 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=131490 $D=0
M1242 378 62 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=126860 $D=0
M1243 379 62 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=131490 $D=0
M1244 6 63 380 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=126860 $D=0
M1245 6 63 381 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=131490 $D=0
M1246 382 64 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=126860 $D=0
M1247 383 64 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=131490 $D=0
M1248 384 380 214 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=126860 $D=0
M1249 385 381 215 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=131490 $D=0
M1250 6 384 720 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=126860 $D=0
M1251 6 385 721 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=131490 $D=0
M1252 386 720 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=126860 $D=0
M1253 387 721 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=131490 $D=0
M1254 384 63 386 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=126860 $D=0
M1255 385 63 387 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=131490 $D=0
M1256 386 382 224 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=126860 $D=0
M1257 387 383 225 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=131490 $D=0
M1258 228 388 386 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=126860 $D=0
M1259 229 389 387 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=131490 $D=0
M1260 388 65 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=126860 $D=0
M1261 389 65 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=131490 $D=0
M1262 6 66 390 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=126860 $D=0
M1263 6 66 391 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=131490 $D=0
M1264 392 67 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=126860 $D=0
M1265 393 67 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=131490 $D=0
M1266 394 390 214 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=126860 $D=0
M1267 395 391 215 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=131490 $D=0
M1268 6 394 722 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=126860 $D=0
M1269 6 395 723 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=131490 $D=0
M1270 396 722 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=126860 $D=0
M1271 397 723 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=131490 $D=0
M1272 394 66 396 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=126860 $D=0
M1273 395 66 397 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=131490 $D=0
M1274 396 392 224 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=126860 $D=0
M1275 397 393 225 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=131490 $D=0
M1276 228 398 396 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=126860 $D=0
M1277 229 399 397 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=131490 $D=0
M1278 398 68 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=126860 $D=0
M1279 399 68 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=131490 $D=0
M1280 6 69 400 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=126860 $D=0
M1281 6 69 401 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=131490 $D=0
M1282 402 70 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=126860 $D=0
M1283 403 70 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=131490 $D=0
M1284 404 400 214 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=126860 $D=0
M1285 405 401 215 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=131490 $D=0
M1286 6 404 724 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=126860 $D=0
M1287 6 405 725 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=131490 $D=0
M1288 406 724 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=126860 $D=0
M1289 407 725 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=131490 $D=0
M1290 404 69 406 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=126860 $D=0
M1291 405 69 407 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=131490 $D=0
M1292 406 402 224 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=126860 $D=0
M1293 407 403 225 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=131490 $D=0
M1294 228 408 406 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=126860 $D=0
M1295 229 409 407 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=131490 $D=0
M1296 408 71 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=126860 $D=0
M1297 409 71 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=131490 $D=0
M1298 6 72 410 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=126860 $D=0
M1299 6 72 411 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=131490 $D=0
M1300 412 73 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=126860 $D=0
M1301 413 73 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=131490 $D=0
M1302 414 410 214 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=126860 $D=0
M1303 415 411 215 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=131490 $D=0
M1304 6 414 726 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=126860 $D=0
M1305 6 415 727 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=131490 $D=0
M1306 416 726 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=126860 $D=0
M1307 417 727 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=131490 $D=0
M1308 414 72 416 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=126860 $D=0
M1309 415 72 417 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=131490 $D=0
M1310 416 412 224 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=126860 $D=0
M1311 417 413 225 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=131490 $D=0
M1312 228 418 416 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=126860 $D=0
M1313 229 419 417 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=131490 $D=0
M1314 418 74 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=126860 $D=0
M1315 419 74 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=131490 $D=0
M1316 6 75 420 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=126860 $D=0
M1317 6 75 421 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=131490 $D=0
M1318 422 76 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=126860 $D=0
M1319 423 76 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=131490 $D=0
M1320 424 420 214 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=126860 $D=0
M1321 425 421 215 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=131490 $D=0
M1322 6 424 728 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=126860 $D=0
M1323 6 425 729 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=131490 $D=0
M1324 426 728 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=126860 $D=0
M1325 427 729 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=131490 $D=0
M1326 424 75 426 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=126860 $D=0
M1327 425 75 427 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=131490 $D=0
M1328 426 422 224 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=126860 $D=0
M1329 427 423 225 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=131490 $D=0
M1330 228 428 426 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=126860 $D=0
M1331 229 429 427 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=131490 $D=0
M1332 428 77 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=126860 $D=0
M1333 429 77 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=131490 $D=0
M1334 6 78 430 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=126860 $D=0
M1335 6 78 431 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=131490 $D=0
M1336 432 79 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=126860 $D=0
M1337 433 79 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=131490 $D=0
M1338 434 430 214 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=126860 $D=0
M1339 435 431 215 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=131490 $D=0
M1340 6 434 730 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=126860 $D=0
M1341 6 435 731 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=131490 $D=0
M1342 436 730 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=126860 $D=0
M1343 437 731 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=131490 $D=0
M1344 434 78 436 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=126860 $D=0
M1345 435 78 437 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=131490 $D=0
M1346 436 432 224 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=126860 $D=0
M1347 437 433 225 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=131490 $D=0
M1348 228 438 436 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=126860 $D=0
M1349 229 439 437 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=131490 $D=0
M1350 438 80 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=126860 $D=0
M1351 439 80 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=131490 $D=0
M1352 6 81 440 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=126860 $D=0
M1353 6 81 441 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=131490 $D=0
M1354 442 82 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=126860 $D=0
M1355 443 82 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=131490 $D=0
M1356 444 440 214 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=126860 $D=0
M1357 445 441 215 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=131490 $D=0
M1358 6 444 732 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=126860 $D=0
M1359 6 445 733 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=131490 $D=0
M1360 446 732 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=126860 $D=0
M1361 447 733 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=131490 $D=0
M1362 444 81 446 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=126860 $D=0
M1363 445 81 447 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=131490 $D=0
M1364 446 442 224 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=126860 $D=0
M1365 447 443 225 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=131490 $D=0
M1366 228 448 446 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=126860 $D=0
M1367 229 449 447 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=131490 $D=0
M1368 448 83 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=126860 $D=0
M1369 449 83 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=131490 $D=0
M1370 6 84 450 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=126860 $D=0
M1371 6 84 451 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=131490 $D=0
M1372 452 85 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=126860 $D=0
M1373 453 85 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=131490 $D=0
M1374 454 450 214 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=126860 $D=0
M1375 455 451 215 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=131490 $D=0
M1376 6 454 734 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=126860 $D=0
M1377 6 455 735 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=131490 $D=0
M1378 456 734 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=126860 $D=0
M1379 457 735 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=131490 $D=0
M1380 454 84 456 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=126860 $D=0
M1381 455 84 457 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=131490 $D=0
M1382 456 452 224 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=126860 $D=0
M1383 457 453 225 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=131490 $D=0
M1384 228 458 456 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=126860 $D=0
M1385 229 459 457 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=131490 $D=0
M1386 458 86 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=126860 $D=0
M1387 459 86 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=131490 $D=0
M1388 6 87 460 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=126860 $D=0
M1389 6 87 461 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=131490 $D=0
M1390 462 88 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=126860 $D=0
M1391 463 88 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=131490 $D=0
M1392 464 460 214 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=126860 $D=0
M1393 465 461 215 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=131490 $D=0
M1394 6 464 736 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=126860 $D=0
M1395 6 465 737 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=131490 $D=0
M1396 466 736 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=126860 $D=0
M1397 467 737 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=131490 $D=0
M1398 464 87 466 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=126860 $D=0
M1399 465 87 467 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=131490 $D=0
M1400 466 462 224 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=126860 $D=0
M1401 467 463 225 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=131490 $D=0
M1402 228 468 466 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=126860 $D=0
M1403 229 469 467 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=131490 $D=0
M1404 468 89 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=126860 $D=0
M1405 469 89 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=131490 $D=0
M1406 6 90 470 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=126860 $D=0
M1407 6 90 471 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=131490 $D=0
M1408 472 91 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=126860 $D=0
M1409 473 91 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=131490 $D=0
M1410 474 470 214 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=126860 $D=0
M1411 475 471 215 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=131490 $D=0
M1412 6 474 738 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=126860 $D=0
M1413 6 475 739 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=131490 $D=0
M1414 476 738 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=126860 $D=0
M1415 477 739 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=131490 $D=0
M1416 474 90 476 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=126860 $D=0
M1417 475 90 477 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=131490 $D=0
M1418 476 472 224 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=126860 $D=0
M1419 477 473 225 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=131490 $D=0
M1420 228 478 476 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=126860 $D=0
M1421 229 479 477 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=131490 $D=0
M1422 478 92 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=126860 $D=0
M1423 479 92 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=131490 $D=0
M1424 6 93 480 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=126860 $D=0
M1425 6 93 481 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=131490 $D=0
M1426 482 94 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=126860 $D=0
M1427 483 94 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=131490 $D=0
M1428 484 480 214 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=126860 $D=0
M1429 485 481 215 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=131490 $D=0
M1430 6 484 740 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=126860 $D=0
M1431 6 485 741 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=131490 $D=0
M1432 486 740 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=126860 $D=0
M1433 487 741 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=131490 $D=0
M1434 484 93 486 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=126860 $D=0
M1435 485 93 487 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=131490 $D=0
M1436 486 482 224 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=126860 $D=0
M1437 487 483 225 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=131490 $D=0
M1438 228 488 486 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=126860 $D=0
M1439 229 489 487 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=131490 $D=0
M1440 488 95 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=126860 $D=0
M1441 489 95 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=131490 $D=0
M1442 6 96 490 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=126860 $D=0
M1443 6 96 491 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=131490 $D=0
M1444 492 97 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=126860 $D=0
M1445 493 97 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=131490 $D=0
M1446 494 490 214 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=126860 $D=0
M1447 495 491 215 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=131490 $D=0
M1448 6 494 742 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=126860 $D=0
M1449 6 495 743 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=131490 $D=0
M1450 496 742 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=126860 $D=0
M1451 497 743 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=131490 $D=0
M1452 494 96 496 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=126860 $D=0
M1453 495 96 497 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=131490 $D=0
M1454 496 492 224 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=126860 $D=0
M1455 497 493 225 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=131490 $D=0
M1456 228 498 496 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=126860 $D=0
M1457 229 499 497 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=131490 $D=0
M1458 498 98 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=126860 $D=0
M1459 499 98 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=131490 $D=0
M1460 6 99 500 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=126860 $D=0
M1461 6 99 501 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=131490 $D=0
M1462 502 100 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=126860 $D=0
M1463 503 100 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=131490 $D=0
M1464 504 500 214 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=126860 $D=0
M1465 505 501 215 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=131490 $D=0
M1466 6 504 744 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=126860 $D=0
M1467 6 505 745 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=131490 $D=0
M1468 506 744 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=126860 $D=0
M1469 507 745 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=131490 $D=0
M1470 504 99 506 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=126860 $D=0
M1471 505 99 507 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=131490 $D=0
M1472 506 502 224 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=126860 $D=0
M1473 507 503 225 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=131490 $D=0
M1474 228 508 506 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=126860 $D=0
M1475 229 509 507 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=131490 $D=0
M1476 508 101 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=126860 $D=0
M1477 509 101 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=131490 $D=0
M1478 6 102 510 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=126860 $D=0
M1479 6 102 511 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=131490 $D=0
M1480 512 103 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=126860 $D=0
M1481 513 103 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=131490 $D=0
M1482 514 510 214 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=126860 $D=0
M1483 515 511 215 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=131490 $D=0
M1484 6 514 746 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=126860 $D=0
M1485 6 515 747 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=131490 $D=0
M1486 516 746 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=126860 $D=0
M1487 517 747 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=131490 $D=0
M1488 514 102 516 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=126860 $D=0
M1489 515 102 517 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=131490 $D=0
M1490 516 512 224 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=126860 $D=0
M1491 517 513 225 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=131490 $D=0
M1492 228 518 516 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=126860 $D=0
M1493 229 519 517 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=131490 $D=0
M1494 518 104 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=126860 $D=0
M1495 519 104 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=131490 $D=0
M1496 6 105 520 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=126860 $D=0
M1497 6 105 521 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=131490 $D=0
M1498 522 106 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=126860 $D=0
M1499 523 106 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=131490 $D=0
M1500 524 520 214 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=126860 $D=0
M1501 525 521 215 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=131490 $D=0
M1502 6 524 748 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=126860 $D=0
M1503 6 525 749 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=131490 $D=0
M1504 526 748 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=126860 $D=0
M1505 527 749 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=131490 $D=0
M1506 524 105 526 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=126860 $D=0
M1507 525 105 527 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=131490 $D=0
M1508 526 522 224 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=126860 $D=0
M1509 527 523 225 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=131490 $D=0
M1510 228 528 526 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=126860 $D=0
M1511 229 529 527 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=131490 $D=0
M1512 528 107 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=126860 $D=0
M1513 529 107 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=131490 $D=0
M1514 6 108 530 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=126860 $D=0
M1515 6 108 531 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=131490 $D=0
M1516 532 109 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=126860 $D=0
M1517 533 109 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=131490 $D=0
M1518 8 532 224 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=126860 $D=0
M1519 8 533 225 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=131490 $D=0
M1520 228 530 8 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=126860 $D=0
M1521 229 531 8 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=131490 $D=0
M1522 6 536 534 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=126860 $D=0
M1523 6 537 535 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=131490 $D=0
M1524 536 110 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=126860 $D=0
M1525 537 110 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=131490 $D=0
M1526 750 224 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=126860 $D=0
M1527 751 225 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=131490 $D=0
M1528 538 536 750 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=126860 $D=0
M1529 539 537 751 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=131490 $D=0
M1530 6 538 540 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=126860 $D=0
M1531 6 539 541 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=131490 $D=0
M1532 752 540 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=126860 $D=0
M1533 753 541 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=131490 $D=0
M1534 538 534 752 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=126860 $D=0
M1535 539 535 753 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=131490 $D=0
M1536 6 544 542 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=126860 $D=0
M1537 6 545 543 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=131490 $D=0
M1538 544 110 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=126860 $D=0
M1539 545 110 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=131490 $D=0
M1540 754 228 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=126860 $D=0
M1541 755 229 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=131490 $D=0
M1542 546 544 754 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=126860 $D=0
M1543 547 545 755 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=131490 $D=0
M1544 6 546 111 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=126860 $D=0
M1545 6 547 112 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=131490 $D=0
M1546 756 111 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=126860 $D=0
M1547 757 112 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=131490 $D=0
M1548 546 542 756 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=126860 $D=0
M1549 547 543 757 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=131490 $D=0
M1550 548 113 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=126860 $D=0
M1551 549 113 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=131490 $D=0
M1552 550 113 540 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=126860 $D=0
M1553 551 113 541 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=131490 $D=0
M1554 114 548 550 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=126860 $D=0
M1555 115 549 551 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=131490 $D=0
M1556 552 116 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=126860 $D=0
M1557 553 116 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=131490 $D=0
M1558 554 116 111 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=126860 $D=0
M1559 555 116 112 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=131490 $D=0
M1560 758 552 554 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=126860 $D=0
M1561 759 553 555 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=131490 $D=0
M1562 6 111 758 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=126860 $D=0
M1563 6 112 759 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=131490 $D=0
M1564 556 117 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=126860 $D=0
M1565 557 117 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=131490 $D=0
M1566 118 117 554 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=126860 $D=0
M1567 119 117 555 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=131490 $D=0
M1568 9 556 118 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=126860 $D=0
M1569 10 557 119 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=131490 $D=0
M1570 559 558 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=126860 $D=0
M1571 560 120 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=131490 $D=0
M1572 6 563 561 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=126860 $D=0
M1573 6 564 562 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=131490 $D=0
M1574 565 550 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=126860 $D=0
M1575 566 551 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=131490 $D=0
M1576 563 550 558 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=126860 $D=0
M1577 564 551 120 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=131490 $D=0
M1578 559 565 563 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=126860 $D=0
M1579 560 566 564 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=131490 $D=0
M1580 567 561 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=126860 $D=0
M1581 568 562 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=131490 $D=0
M1582 121 561 118 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=126860 $D=0
M1583 558 562 119 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=131490 $D=0
M1584 550 567 121 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=126860 $D=0
M1585 551 568 558 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=131490 $D=0
M1586 569 121 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=126860 $D=0
M1587 570 558 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=131490 $D=0
M1588 571 561 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=126860 $D=0
M1589 572 562 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=131490 $D=0
M1590 573 561 569 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=126860 $D=0
M1591 574 562 570 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=131490 $D=0
M1592 118 571 573 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=126860 $D=0
M1593 119 572 574 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=131490 $D=0
M1594 770 550 6 6 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=126500 $D=0
M1595 771 551 6 6 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=131130 $D=0
M1596 575 118 770 6 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=126500 $D=0
M1597 576 119 771 6 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=131130 $D=0
M1598 577 573 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=126860 $D=0
M1599 578 574 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=131490 $D=0
M1600 579 550 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=126860 $D=0
M1601 580 551 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=131490 $D=0
M1602 6 118 579 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=126860 $D=0
M1603 6 119 580 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=131490 $D=0
M1604 581 550 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=126860 $D=0
M1605 582 551 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=131490 $D=0
M1606 6 118 581 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=126860 $D=0
M1607 6 119 582 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=131490 $D=0
M1608 772 550 6 6 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=126680 $D=0
M1609 773 551 6 6 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=131310 $D=0
M1610 585 118 772 6 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=126680 $D=0
M1611 586 119 773 6 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=131310 $D=0
M1612 6 581 585 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=126860 $D=0
M1613 6 582 586 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=131490 $D=0
M1614 587 127 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=126860 $D=0
M1615 588 127 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=131490 $D=0
M1616 589 127 575 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=126860 $D=0
M1617 590 127 576 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=131490 $D=0
M1618 579 587 589 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=126860 $D=0
M1619 580 588 590 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=131490 $D=0
M1620 591 127 577 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=126860 $D=0
M1621 592 127 578 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=131490 $D=0
M1622 585 587 591 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=126860 $D=0
M1623 586 588 592 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=131490 $D=0
M1624 593 128 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=126860 $D=0
M1625 594 128 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=131490 $D=0
M1626 595 128 591 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=126860 $D=0
M1627 596 128 592 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=131490 $D=0
M1628 589 593 595 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=126860 $D=0
M1629 590 594 596 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=131490 $D=0
M1630 11 595 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=126860 $D=0
M1631 12 596 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=131490 $D=0
M1632 597 130 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=126860 $D=0
M1633 598 130 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=131490 $D=0
M1634 599 130 131 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=126860 $D=0
M1635 600 130 132 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=131490 $D=0
M1636 133 597 599 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=126860 $D=0
M1637 134 598 600 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=131490 $D=0
M1638 601 130 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=126860 $D=0
M1639 602 130 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=131490 $D=0
M1640 603 130 135 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=126860 $D=0
M1641 604 130 136 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=131490 $D=0
M1642 137 601 603 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=126860 $D=0
M1643 138 602 604 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=131490 $D=0
M1644 605 130 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=126860 $D=0
M1645 606 130 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=131490 $D=0
M1646 607 130 124 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=126860 $D=0
M1647 608 130 8 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=131490 $D=0
M1648 129 605 607 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=126860 $D=0
M1649 139 606 608 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=131490 $D=0
M1650 609 130 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=126860 $D=0
M1651 610 130 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=131490 $D=0
M1652 611 130 8 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=126860 $D=0
M1653 612 130 8 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=131490 $D=0
M1654 140 609 611 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=126860 $D=0
M1655 141 610 612 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=131490 $D=0
M1656 613 130 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=126860 $D=0
M1657 614 130 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=131490 $D=0
M1658 615 130 8 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=126860 $D=0
M1659 616 130 8 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=131490 $D=0
M1660 142 613 615 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=126860 $D=0
M1661 143 614 616 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=131490 $D=0
M1662 6 550 760 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=126860 $D=0
M1663 6 551 761 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=131490 $D=0
M1664 134 760 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=126860 $D=0
M1665 131 761 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=131490 $D=0
M1666 617 144 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=126860 $D=0
M1667 618 144 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=131490 $D=0
M1668 145 144 134 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=126860 $D=0
M1669 146 144 131 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=131490 $D=0
M1670 599 617 145 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=126860 $D=0
M1671 600 618 146 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=131490 $D=0
M1672 619 147 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=126860 $D=0
M1673 620 147 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=131490 $D=0
M1674 148 147 145 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=126860 $D=0
M1675 126 147 146 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=131490 $D=0
M1676 603 619 148 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=126860 $D=0
M1677 604 620 126 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=131490 $D=0
M1678 621 149 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=126860 $D=0
M1679 622 149 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=131490 $D=0
M1680 122 149 148 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=126860 $D=0
M1681 123 149 126 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=131490 $D=0
M1682 607 621 122 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=126860 $D=0
M1683 608 622 123 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=131490 $D=0
M1684 623 119 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=126860 $D=0
M1685 624 119 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=131490 $D=0
M1686 150 119 122 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=126860 $D=0
M1687 151 119 123 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=131490 $D=0
M1688 611 623 150 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=126860 $D=0
M1689 612 624 151 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=131490 $D=0
M1690 625 118 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=126860 $D=0
M1691 626 118 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=131490 $D=0
M1692 200 118 150 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=126860 $D=0
M1693 201 118 151 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=131490 $D=0
M1694 615 625 200 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=126860 $D=0
M1695 616 626 201 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=131490 $D=0
M1696 627 152 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=126860 $D=0
M1697 628 152 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=131490 $D=0
M1698 629 152 111 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=126860 $D=0
M1699 630 152 112 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=131490 $D=0
M1700 9 627 629 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=126860 $D=0
M1701 10 628 630 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=131490 $D=0
M1702 631 540 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=126860 $D=0
M1703 632 541 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=131490 $D=0
M1704 6 629 631 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=126860 $D=0
M1705 6 630 632 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=131490 $D=0
M1706 774 540 6 6 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=126680 $D=0
M1707 775 541 6 6 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=131310 $D=0
M1708 635 629 774 6 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=126680 $D=0
M1709 636 630 775 6 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=131310 $D=0
M1710 6 631 635 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=126860 $D=0
M1711 6 632 636 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=131490 $D=0
M1712 762 153 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=126860 $D=0
M1713 763 637 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=131490 $D=0
M1714 6 635 762 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=126860 $D=0
M1715 6 636 763 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=131490 $D=0
M1716 637 762 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=126860 $D=0
M1717 154 763 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=131490 $D=0
M1718 776 540 6 6 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=126500 $D=0
M1719 777 541 6 6 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=131130 $D=0
M1720 638 640 776 6 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=126500 $D=0
M1721 639 641 777 6 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=131130 $D=0
M1722 640 629 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=126860 $D=0
M1723 641 630 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=131490 $D=0
M1724 642 638 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=126860 $D=0
M1725 643 639 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=131490 $D=0
M1726 6 153 642 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=126860 $D=0
M1727 6 637 643 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=131490 $D=0
M1728 645 155 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=126860 $D=0
M1729 646 644 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=131490 $D=0
M1730 644 642 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=126860 $D=0
M1731 156 643 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=131490 $D=0
M1732 6 645 644 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=126860 $D=0
M1733 6 646 156 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=131490 $D=0
M1734 648 647 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=126860 $D=0
M1735 649 157 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=131490 $D=0
M1736 6 652 650 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=126860 $D=0
M1737 6 653 651 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=131490 $D=0
M1738 654 114 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=126860 $D=0
M1739 655 115 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=131490 $D=0
M1740 652 114 647 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=126860 $D=0
M1741 653 115 157 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=131490 $D=0
M1742 648 654 652 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=126860 $D=0
M1743 649 655 653 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=131490 $D=0
M1744 656 650 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=126860 $D=0
M1745 657 651 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=131490 $D=0
M1746 158 650 8 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=126860 $D=0
M1747 647 651 8 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=131490 $D=0
M1748 114 656 158 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=126860 $D=0
M1749 115 657 647 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=131490 $D=0
M1750 658 158 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=126860 $D=0
M1751 659 647 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=131490 $D=0
M1752 660 650 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=126860 $D=0
M1753 661 651 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=131490 $D=0
M1754 202 650 658 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=126860 $D=0
M1755 203 651 659 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=131490 $D=0
M1756 8 660 202 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=126860 $D=0
M1757 8 661 203 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=131490 $D=0
M1758 662 159 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=126860 $D=0
M1759 663 159 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=131490 $D=0
M1760 664 159 202 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=126860 $D=0
M1761 665 159 203 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=131490 $D=0
M1762 11 662 664 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=126860 $D=0
M1763 12 663 665 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=131490 $D=0
M1764 666 160 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=126860 $D=0
M1765 667 160 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=131490 $D=0
M1766 668 160 664 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=126860 $D=0
M1767 669 160 665 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=131490 $D=0
M1768 8 666 668 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=126860 $D=0
M1769 8 667 669 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=131490 $D=0
M1770 670 110 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=126860 $D=0
M1771 671 110 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=131490 $D=0
M1772 6 670 672 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=126860 $D=0
M1773 6 671 673 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=131490 $D=0
M1774 674 110 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=126860 $D=0
M1775 675 110 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=131490 $D=0
M1776 676 672 668 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=126860 $D=0
M1777 677 673 669 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=131490 $D=0
M1778 6 676 764 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=126860 $D=0
M1779 6 677 765 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=131490 $D=0
M1780 678 764 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=126860 $D=0
M1781 679 765 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=131490 $D=0
M1782 676 670 678 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=126860 $D=0
M1783 677 671 679 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=131490 $D=0
M1784 680 674 678 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=126860 $D=0
M1785 681 675 679 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=131490 $D=0
M1786 6 684 682 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=126860 $D=0
M1787 6 685 683 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=131490 $D=0
M1788 684 110 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=126860 $D=0
M1789 685 110 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=131490 $D=0
M1790 766 680 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=126860 $D=0
M1791 767 681 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=131490 $D=0
M1792 686 684 766 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=126860 $D=0
M1793 687 685 767 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=131490 $D=0
M1794 6 686 114 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=126860 $D=0
M1795 6 687 115 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=131490 $D=0
M1796 768 114 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=126860 $D=0
M1797 769 115 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=131490 $D=0
M1798 686 682 768 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=126860 $D=0
M1799 687 683 769 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=131490 $D=0
.ENDS
***************************************
.SUBCKT ICV_26 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141
+ 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161
** N=800 EP=160 IP=1514 FDC=1800
M0 185 1 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=116350 $D=1
M1 186 1 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=120980 $D=1
M2 187 185 2 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=116350 $D=1
M3 188 186 3 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=120980 $D=1
M4 8 1 187 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=116350 $D=1
M5 8 1 188 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=120980 $D=1
M6 189 185 2 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=116350 $D=1
M7 190 186 3 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=120980 $D=1
M8 2 1 189 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=116350 $D=1
M9 3 1 190 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=120980 $D=1
M10 191 185 2 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=116350 $D=1
M11 192 186 3 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=120980 $D=1
M12 2 1 191 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=116350 $D=1
M13 3 1 192 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=120980 $D=1
M14 195 193 191 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=116350 $D=1
M15 196 194 192 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=120980 $D=1
M16 193 4 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=116350 $D=1
M17 194 4 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=120980 $D=1
M18 197 193 189 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=116350 $D=1
M19 198 194 190 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=120980 $D=1
M20 187 4 197 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=116350 $D=1
M21 188 4 198 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=120980 $D=1
M22 199 5 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=116350 $D=1
M23 200 5 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=120980 $D=1
M24 201 199 197 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=116350 $D=1
M25 202 200 198 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=120980 $D=1
M26 195 5 201 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=116350 $D=1
M27 196 5 202 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=120980 $D=1
M28 203 7 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=116350 $D=1
M29 204 7 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=120980 $D=1
M30 205 203 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=116350 $D=1
M31 206 204 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=120980 $D=1
M32 9 7 205 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=116350 $D=1
M33 10 7 206 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=120980 $D=1
M34 207 203 11 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=116350 $D=1
M35 208 204 12 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=120980 $D=1
M36 209 7 207 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=116350 $D=1
M37 210 7 208 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=120980 $D=1
M38 213 203 211 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=116350 $D=1
M39 214 204 212 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=120980 $D=1
M40 201 7 213 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=116350 $D=1
M41 202 7 214 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=120980 $D=1
M42 217 215 213 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=116350 $D=1
M43 218 216 214 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=120980 $D=1
M44 215 13 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=116350 $D=1
M45 216 13 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=120980 $D=1
M46 219 215 207 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=116350 $D=1
M47 220 216 208 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=120980 $D=1
M48 205 13 219 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=116350 $D=1
M49 206 13 220 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=120980 $D=1
M50 221 14 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=116350 $D=1
M51 222 14 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=120980 $D=1
M52 223 221 219 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=116350 $D=1
M53 224 222 220 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=120980 $D=1
M54 217 14 223 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=116350 $D=1
M55 218 14 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=120980 $D=1
M56 8 15 225 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=116350 $D=1
M57 8 15 226 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=120980 $D=1
M58 227 16 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=116350 $D=1
M59 228 16 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=120980 $D=1
M60 229 15 223 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=116350 $D=1
M61 230 15 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=120980 $D=1
M62 8 229 699 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=116350 $D=1
M63 8 230 700 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=120980 $D=1
M64 231 699 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=116350 $D=1
M65 232 700 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=120980 $D=1
M66 229 225 231 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=116350 $D=1
M67 230 226 232 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=120980 $D=1
M68 231 16 233 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=116350 $D=1
M69 232 16 234 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=120980 $D=1
M70 237 17 231 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=116350 $D=1
M71 238 17 232 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=120980 $D=1
M72 235 17 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=116350 $D=1
M73 236 17 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=120980 $D=1
M74 8 18 239 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=116350 $D=1
M75 8 18 240 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=120980 $D=1
M76 241 19 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=116350 $D=1
M77 242 19 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=120980 $D=1
M78 243 18 223 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=116350 $D=1
M79 244 18 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=120980 $D=1
M80 8 243 701 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=116350 $D=1
M81 8 244 702 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=120980 $D=1
M82 245 701 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=116350 $D=1
M83 246 702 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=120980 $D=1
M84 243 239 245 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=116350 $D=1
M85 244 240 246 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=120980 $D=1
M86 245 19 233 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=116350 $D=1
M87 246 19 234 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=120980 $D=1
M88 237 20 245 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=116350 $D=1
M89 238 20 246 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=120980 $D=1
M90 247 20 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=116350 $D=1
M91 248 20 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=120980 $D=1
M92 8 21 249 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=116350 $D=1
M93 8 21 250 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=120980 $D=1
M94 251 22 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=116350 $D=1
M95 252 22 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=120980 $D=1
M96 253 21 223 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=116350 $D=1
M97 254 21 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=120980 $D=1
M98 8 253 703 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=116350 $D=1
M99 8 254 704 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=120980 $D=1
M100 255 703 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=116350 $D=1
M101 256 704 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=120980 $D=1
M102 253 249 255 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=116350 $D=1
M103 254 250 256 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=120980 $D=1
M104 255 22 233 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=116350 $D=1
M105 256 22 234 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=120980 $D=1
M106 237 23 255 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=116350 $D=1
M107 238 23 256 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=120980 $D=1
M108 257 23 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=116350 $D=1
M109 258 23 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=120980 $D=1
M110 8 24 259 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=116350 $D=1
M111 8 24 260 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=120980 $D=1
M112 261 25 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=116350 $D=1
M113 262 25 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=120980 $D=1
M114 263 24 223 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=116350 $D=1
M115 264 24 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=120980 $D=1
M116 8 263 705 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=116350 $D=1
M117 8 264 706 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=120980 $D=1
M118 265 705 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=116350 $D=1
M119 266 706 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=120980 $D=1
M120 263 259 265 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=116350 $D=1
M121 264 260 266 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=120980 $D=1
M122 265 25 233 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=116350 $D=1
M123 266 25 234 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=120980 $D=1
M124 237 26 265 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=116350 $D=1
M125 238 26 266 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=120980 $D=1
M126 267 26 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=116350 $D=1
M127 268 26 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=120980 $D=1
M128 8 27 269 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=116350 $D=1
M129 8 27 270 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=120980 $D=1
M130 271 28 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=116350 $D=1
M131 272 28 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=120980 $D=1
M132 273 27 223 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=116350 $D=1
M133 274 27 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=120980 $D=1
M134 8 273 707 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=116350 $D=1
M135 8 274 708 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=120980 $D=1
M136 275 707 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=116350 $D=1
M137 276 708 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=120980 $D=1
M138 273 269 275 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=116350 $D=1
M139 274 270 276 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=120980 $D=1
M140 275 28 233 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=116350 $D=1
M141 276 28 234 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=120980 $D=1
M142 237 29 275 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=116350 $D=1
M143 238 29 276 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=120980 $D=1
M144 277 29 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=116350 $D=1
M145 278 29 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=120980 $D=1
M146 8 30 279 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=116350 $D=1
M147 8 30 280 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=120980 $D=1
M148 281 31 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=116350 $D=1
M149 282 31 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=120980 $D=1
M150 283 30 223 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=116350 $D=1
M151 284 30 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=120980 $D=1
M152 8 283 709 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=116350 $D=1
M153 8 284 710 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=120980 $D=1
M154 285 709 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=116350 $D=1
M155 286 710 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=120980 $D=1
M156 283 279 285 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=116350 $D=1
M157 284 280 286 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=120980 $D=1
M158 285 31 233 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=116350 $D=1
M159 286 31 234 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=120980 $D=1
M160 237 32 285 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=116350 $D=1
M161 238 32 286 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=120980 $D=1
M162 287 32 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=116350 $D=1
M163 288 32 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=120980 $D=1
M164 8 33 289 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=116350 $D=1
M165 8 33 290 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=120980 $D=1
M166 291 34 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=116350 $D=1
M167 292 34 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=120980 $D=1
M168 293 33 223 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=116350 $D=1
M169 294 33 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=120980 $D=1
M170 8 293 711 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=116350 $D=1
M171 8 294 712 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=120980 $D=1
M172 295 711 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=116350 $D=1
M173 296 712 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=120980 $D=1
M174 293 289 295 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=116350 $D=1
M175 294 290 296 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=120980 $D=1
M176 295 34 233 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=116350 $D=1
M177 296 34 234 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=120980 $D=1
M178 237 35 295 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=116350 $D=1
M179 238 35 296 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=120980 $D=1
M180 297 35 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=116350 $D=1
M181 298 35 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=120980 $D=1
M182 8 36 299 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=116350 $D=1
M183 8 36 300 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=120980 $D=1
M184 301 37 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=116350 $D=1
M185 302 37 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=120980 $D=1
M186 303 36 223 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=116350 $D=1
M187 304 36 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=120980 $D=1
M188 8 303 713 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=116350 $D=1
M189 8 304 714 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=120980 $D=1
M190 305 713 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=116350 $D=1
M191 306 714 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=120980 $D=1
M192 303 299 305 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=116350 $D=1
M193 304 300 306 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=120980 $D=1
M194 305 37 233 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=116350 $D=1
M195 306 37 234 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=120980 $D=1
M196 237 38 305 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=116350 $D=1
M197 238 38 306 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=120980 $D=1
M198 307 38 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=116350 $D=1
M199 308 38 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=120980 $D=1
M200 8 39 309 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=116350 $D=1
M201 8 39 310 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=120980 $D=1
M202 311 40 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=116350 $D=1
M203 312 40 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=120980 $D=1
M204 313 39 223 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=116350 $D=1
M205 314 39 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=120980 $D=1
M206 8 313 715 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=116350 $D=1
M207 8 314 716 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=120980 $D=1
M208 315 715 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=116350 $D=1
M209 316 716 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=120980 $D=1
M210 313 309 315 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=116350 $D=1
M211 314 310 316 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=120980 $D=1
M212 315 40 233 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=116350 $D=1
M213 316 40 234 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=120980 $D=1
M214 237 41 315 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=116350 $D=1
M215 238 41 316 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=120980 $D=1
M216 317 41 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=116350 $D=1
M217 318 41 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=120980 $D=1
M218 8 42 319 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=116350 $D=1
M219 8 42 320 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=120980 $D=1
M220 321 43 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=116350 $D=1
M221 322 43 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=120980 $D=1
M222 323 42 223 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=116350 $D=1
M223 324 42 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=120980 $D=1
M224 8 323 717 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=116350 $D=1
M225 8 324 718 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=120980 $D=1
M226 325 717 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=116350 $D=1
M227 326 718 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=120980 $D=1
M228 323 319 325 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=116350 $D=1
M229 324 320 326 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=120980 $D=1
M230 325 43 233 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=116350 $D=1
M231 326 43 234 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=120980 $D=1
M232 237 44 325 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=116350 $D=1
M233 238 44 326 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=120980 $D=1
M234 327 44 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=116350 $D=1
M235 328 44 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=120980 $D=1
M236 8 45 329 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=116350 $D=1
M237 8 45 330 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=120980 $D=1
M238 331 46 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=116350 $D=1
M239 332 46 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=120980 $D=1
M240 333 45 223 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=116350 $D=1
M241 334 45 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=120980 $D=1
M242 8 333 719 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=116350 $D=1
M243 8 334 720 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=120980 $D=1
M244 335 719 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=116350 $D=1
M245 336 720 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=120980 $D=1
M246 333 329 335 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=116350 $D=1
M247 334 330 336 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=120980 $D=1
M248 335 46 233 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=116350 $D=1
M249 336 46 234 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=120980 $D=1
M250 237 47 335 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=116350 $D=1
M251 238 47 336 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=120980 $D=1
M252 337 47 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=116350 $D=1
M253 338 47 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=120980 $D=1
M254 8 48 339 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=116350 $D=1
M255 8 48 340 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=120980 $D=1
M256 341 49 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=116350 $D=1
M257 342 49 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=120980 $D=1
M258 343 48 223 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=116350 $D=1
M259 344 48 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=120980 $D=1
M260 8 343 721 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=116350 $D=1
M261 8 344 722 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=120980 $D=1
M262 345 721 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=116350 $D=1
M263 346 722 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=120980 $D=1
M264 343 339 345 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=116350 $D=1
M265 344 340 346 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=120980 $D=1
M266 345 49 233 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=116350 $D=1
M267 346 49 234 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=120980 $D=1
M268 237 50 345 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=116350 $D=1
M269 238 50 346 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=120980 $D=1
M270 347 50 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=116350 $D=1
M271 348 50 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=120980 $D=1
M272 8 51 349 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=116350 $D=1
M273 8 51 350 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=120980 $D=1
M274 351 52 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=116350 $D=1
M275 352 52 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=120980 $D=1
M276 353 51 223 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=116350 $D=1
M277 354 51 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=120980 $D=1
M278 8 353 723 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=116350 $D=1
M279 8 354 724 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=120980 $D=1
M280 355 723 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=116350 $D=1
M281 356 724 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=120980 $D=1
M282 353 349 355 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=116350 $D=1
M283 354 350 356 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=120980 $D=1
M284 355 52 233 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=116350 $D=1
M285 356 52 234 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=120980 $D=1
M286 237 53 355 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=116350 $D=1
M287 238 53 356 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=120980 $D=1
M288 357 53 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=116350 $D=1
M289 358 53 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=120980 $D=1
M290 8 54 359 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=116350 $D=1
M291 8 54 360 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=120980 $D=1
M292 361 55 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=116350 $D=1
M293 362 55 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=120980 $D=1
M294 363 54 223 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=116350 $D=1
M295 364 54 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=120980 $D=1
M296 8 363 725 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=116350 $D=1
M297 8 364 726 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=120980 $D=1
M298 365 725 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=116350 $D=1
M299 366 726 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=120980 $D=1
M300 363 359 365 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=116350 $D=1
M301 364 360 366 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=120980 $D=1
M302 365 55 233 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=116350 $D=1
M303 366 55 234 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=120980 $D=1
M304 237 56 365 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=116350 $D=1
M305 238 56 366 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=120980 $D=1
M306 367 56 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=116350 $D=1
M307 368 56 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=120980 $D=1
M308 8 57 369 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=116350 $D=1
M309 8 57 370 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=120980 $D=1
M310 371 58 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=116350 $D=1
M311 372 58 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=120980 $D=1
M312 373 57 223 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=116350 $D=1
M313 374 57 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=120980 $D=1
M314 8 373 727 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=116350 $D=1
M315 8 374 728 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=120980 $D=1
M316 375 727 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=116350 $D=1
M317 376 728 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=120980 $D=1
M318 373 369 375 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=116350 $D=1
M319 374 370 376 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=120980 $D=1
M320 375 58 233 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=116350 $D=1
M321 376 58 234 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=120980 $D=1
M322 237 59 375 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=116350 $D=1
M323 238 59 376 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=120980 $D=1
M324 377 59 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=116350 $D=1
M325 378 59 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=120980 $D=1
M326 8 60 379 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=116350 $D=1
M327 8 60 380 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=120980 $D=1
M328 381 61 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=116350 $D=1
M329 382 61 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=120980 $D=1
M330 383 60 223 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=116350 $D=1
M331 384 60 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=120980 $D=1
M332 8 383 729 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=116350 $D=1
M333 8 384 730 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=120980 $D=1
M334 385 729 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=116350 $D=1
M335 386 730 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=120980 $D=1
M336 383 379 385 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=116350 $D=1
M337 384 380 386 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=120980 $D=1
M338 385 61 233 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=116350 $D=1
M339 386 61 234 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=120980 $D=1
M340 237 62 385 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=116350 $D=1
M341 238 62 386 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=120980 $D=1
M342 387 62 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=116350 $D=1
M343 388 62 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=120980 $D=1
M344 8 63 389 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=116350 $D=1
M345 8 63 390 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=120980 $D=1
M346 391 64 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=116350 $D=1
M347 392 64 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=120980 $D=1
M348 393 63 223 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=116350 $D=1
M349 394 63 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=120980 $D=1
M350 8 393 731 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=116350 $D=1
M351 8 394 732 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=120980 $D=1
M352 395 731 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=116350 $D=1
M353 396 732 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=120980 $D=1
M354 393 389 395 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=116350 $D=1
M355 394 390 396 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=120980 $D=1
M356 395 64 233 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=116350 $D=1
M357 396 64 234 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=120980 $D=1
M358 237 65 395 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=116350 $D=1
M359 238 65 396 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=120980 $D=1
M360 397 65 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=116350 $D=1
M361 398 65 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=120980 $D=1
M362 8 66 399 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=116350 $D=1
M363 8 66 400 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=120980 $D=1
M364 401 67 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=116350 $D=1
M365 402 67 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=120980 $D=1
M366 403 66 223 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=116350 $D=1
M367 404 66 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=120980 $D=1
M368 8 403 733 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=116350 $D=1
M369 8 404 734 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=120980 $D=1
M370 405 733 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=116350 $D=1
M371 406 734 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=120980 $D=1
M372 403 399 405 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=116350 $D=1
M373 404 400 406 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=120980 $D=1
M374 405 67 233 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=116350 $D=1
M375 406 67 234 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=120980 $D=1
M376 237 68 405 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=116350 $D=1
M377 238 68 406 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=120980 $D=1
M378 407 68 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=116350 $D=1
M379 408 68 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=120980 $D=1
M380 8 69 409 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=116350 $D=1
M381 8 69 410 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=120980 $D=1
M382 411 70 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=116350 $D=1
M383 412 70 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=120980 $D=1
M384 413 69 223 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=116350 $D=1
M385 414 69 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=120980 $D=1
M386 8 413 735 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=116350 $D=1
M387 8 414 736 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=120980 $D=1
M388 415 735 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=116350 $D=1
M389 416 736 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=120980 $D=1
M390 413 409 415 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=116350 $D=1
M391 414 410 416 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=120980 $D=1
M392 415 70 233 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=116350 $D=1
M393 416 70 234 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=120980 $D=1
M394 237 71 415 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=116350 $D=1
M395 238 71 416 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=120980 $D=1
M396 417 71 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=116350 $D=1
M397 418 71 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=120980 $D=1
M398 8 72 419 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=116350 $D=1
M399 8 72 420 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=120980 $D=1
M400 421 73 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=116350 $D=1
M401 422 73 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=120980 $D=1
M402 423 72 223 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=116350 $D=1
M403 424 72 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=120980 $D=1
M404 8 423 737 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=116350 $D=1
M405 8 424 738 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=120980 $D=1
M406 425 737 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=116350 $D=1
M407 426 738 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=120980 $D=1
M408 423 419 425 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=116350 $D=1
M409 424 420 426 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=120980 $D=1
M410 425 73 233 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=116350 $D=1
M411 426 73 234 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=120980 $D=1
M412 237 74 425 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=116350 $D=1
M413 238 74 426 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=120980 $D=1
M414 427 74 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=116350 $D=1
M415 428 74 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=120980 $D=1
M416 8 75 429 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=116350 $D=1
M417 8 75 430 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=120980 $D=1
M418 431 76 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=116350 $D=1
M419 432 76 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=120980 $D=1
M420 433 75 223 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=116350 $D=1
M421 434 75 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=120980 $D=1
M422 8 433 739 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=116350 $D=1
M423 8 434 740 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=120980 $D=1
M424 435 739 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=116350 $D=1
M425 436 740 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=120980 $D=1
M426 433 429 435 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=116350 $D=1
M427 434 430 436 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=120980 $D=1
M428 435 76 233 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=116350 $D=1
M429 436 76 234 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=120980 $D=1
M430 237 77 435 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=116350 $D=1
M431 238 77 436 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=120980 $D=1
M432 437 77 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=116350 $D=1
M433 438 77 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=120980 $D=1
M434 8 78 439 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=116350 $D=1
M435 8 78 440 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=120980 $D=1
M436 441 79 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=116350 $D=1
M437 442 79 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=120980 $D=1
M438 443 78 223 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=116350 $D=1
M439 444 78 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=120980 $D=1
M440 8 443 741 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=116350 $D=1
M441 8 444 742 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=120980 $D=1
M442 445 741 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=116350 $D=1
M443 446 742 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=120980 $D=1
M444 443 439 445 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=116350 $D=1
M445 444 440 446 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=120980 $D=1
M446 445 79 233 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=116350 $D=1
M447 446 79 234 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=120980 $D=1
M448 237 80 445 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=116350 $D=1
M449 238 80 446 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=120980 $D=1
M450 447 80 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=116350 $D=1
M451 448 80 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=120980 $D=1
M452 8 81 449 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=116350 $D=1
M453 8 81 450 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=120980 $D=1
M454 451 82 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=116350 $D=1
M455 452 82 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=120980 $D=1
M456 453 81 223 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=116350 $D=1
M457 454 81 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=120980 $D=1
M458 8 453 743 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=116350 $D=1
M459 8 454 744 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=120980 $D=1
M460 455 743 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=116350 $D=1
M461 456 744 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=120980 $D=1
M462 453 449 455 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=116350 $D=1
M463 454 450 456 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=120980 $D=1
M464 455 82 233 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=116350 $D=1
M465 456 82 234 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=120980 $D=1
M466 237 83 455 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=116350 $D=1
M467 238 83 456 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=120980 $D=1
M468 457 83 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=116350 $D=1
M469 458 83 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=120980 $D=1
M470 8 84 459 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=116350 $D=1
M471 8 84 460 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=120980 $D=1
M472 461 85 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=116350 $D=1
M473 462 85 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=120980 $D=1
M474 463 84 223 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=116350 $D=1
M475 464 84 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=120980 $D=1
M476 8 463 745 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=116350 $D=1
M477 8 464 746 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=120980 $D=1
M478 465 745 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=116350 $D=1
M479 466 746 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=120980 $D=1
M480 463 459 465 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=116350 $D=1
M481 464 460 466 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=120980 $D=1
M482 465 85 233 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=116350 $D=1
M483 466 85 234 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=120980 $D=1
M484 237 86 465 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=116350 $D=1
M485 238 86 466 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=120980 $D=1
M486 467 86 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=116350 $D=1
M487 468 86 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=120980 $D=1
M488 8 87 469 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=116350 $D=1
M489 8 87 470 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=120980 $D=1
M490 471 88 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=116350 $D=1
M491 472 88 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=120980 $D=1
M492 473 87 223 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=116350 $D=1
M493 474 87 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=120980 $D=1
M494 8 473 747 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=116350 $D=1
M495 8 474 748 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=120980 $D=1
M496 475 747 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=116350 $D=1
M497 476 748 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=120980 $D=1
M498 473 469 475 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=116350 $D=1
M499 474 470 476 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=120980 $D=1
M500 475 88 233 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=116350 $D=1
M501 476 88 234 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=120980 $D=1
M502 237 89 475 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=116350 $D=1
M503 238 89 476 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=120980 $D=1
M504 477 89 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=116350 $D=1
M505 478 89 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=120980 $D=1
M506 8 90 479 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=116350 $D=1
M507 8 90 480 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=120980 $D=1
M508 481 91 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=116350 $D=1
M509 482 91 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=120980 $D=1
M510 483 90 223 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=116350 $D=1
M511 484 90 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=120980 $D=1
M512 8 483 749 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=116350 $D=1
M513 8 484 750 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=120980 $D=1
M514 485 749 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=116350 $D=1
M515 486 750 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=120980 $D=1
M516 483 479 485 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=116350 $D=1
M517 484 480 486 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=120980 $D=1
M518 485 91 233 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=116350 $D=1
M519 486 91 234 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=120980 $D=1
M520 237 92 485 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=116350 $D=1
M521 238 92 486 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=120980 $D=1
M522 487 92 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=116350 $D=1
M523 488 92 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=120980 $D=1
M524 8 93 489 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=116350 $D=1
M525 8 93 490 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=120980 $D=1
M526 491 94 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=116350 $D=1
M527 492 94 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=120980 $D=1
M528 493 93 223 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=116350 $D=1
M529 494 93 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=120980 $D=1
M530 8 493 751 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=116350 $D=1
M531 8 494 752 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=120980 $D=1
M532 495 751 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=116350 $D=1
M533 496 752 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=120980 $D=1
M534 493 489 495 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=116350 $D=1
M535 494 490 496 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=120980 $D=1
M536 495 94 233 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=116350 $D=1
M537 496 94 234 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=120980 $D=1
M538 237 95 495 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=116350 $D=1
M539 238 95 496 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=120980 $D=1
M540 497 95 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=116350 $D=1
M541 498 95 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=120980 $D=1
M542 8 96 499 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=116350 $D=1
M543 8 96 500 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=120980 $D=1
M544 501 97 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=116350 $D=1
M545 502 97 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=120980 $D=1
M546 503 96 223 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=116350 $D=1
M547 504 96 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=120980 $D=1
M548 8 503 753 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=116350 $D=1
M549 8 504 754 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=120980 $D=1
M550 505 753 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=116350 $D=1
M551 506 754 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=120980 $D=1
M552 503 499 505 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=116350 $D=1
M553 504 500 506 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=120980 $D=1
M554 505 97 233 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=116350 $D=1
M555 506 97 234 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=120980 $D=1
M556 237 98 505 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=116350 $D=1
M557 238 98 506 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=120980 $D=1
M558 507 98 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=116350 $D=1
M559 508 98 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=120980 $D=1
M560 8 99 509 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=116350 $D=1
M561 8 99 510 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=120980 $D=1
M562 511 100 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=116350 $D=1
M563 512 100 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=120980 $D=1
M564 513 99 223 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=116350 $D=1
M565 514 99 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=120980 $D=1
M566 8 513 755 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=116350 $D=1
M567 8 514 756 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=120980 $D=1
M568 515 755 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=116350 $D=1
M569 516 756 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=120980 $D=1
M570 513 509 515 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=116350 $D=1
M571 514 510 516 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=120980 $D=1
M572 515 100 233 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=116350 $D=1
M573 516 100 234 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=120980 $D=1
M574 237 101 515 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=116350 $D=1
M575 238 101 516 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=120980 $D=1
M576 517 101 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=116350 $D=1
M577 518 101 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=120980 $D=1
M578 8 102 519 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=116350 $D=1
M579 8 102 520 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=120980 $D=1
M580 521 103 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=116350 $D=1
M581 522 103 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=120980 $D=1
M582 523 102 223 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=116350 $D=1
M583 524 102 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=120980 $D=1
M584 8 523 757 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=116350 $D=1
M585 8 524 758 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=120980 $D=1
M586 525 757 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=116350 $D=1
M587 526 758 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=120980 $D=1
M588 523 519 525 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=116350 $D=1
M589 524 520 526 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=120980 $D=1
M590 525 103 233 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=116350 $D=1
M591 526 103 234 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=120980 $D=1
M592 237 104 525 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=116350 $D=1
M593 238 104 526 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=120980 $D=1
M594 527 104 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=116350 $D=1
M595 528 104 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=120980 $D=1
M596 8 105 529 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=116350 $D=1
M597 8 105 530 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=120980 $D=1
M598 531 106 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=116350 $D=1
M599 532 106 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=120980 $D=1
M600 533 105 223 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=116350 $D=1
M601 534 105 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=120980 $D=1
M602 8 533 759 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=116350 $D=1
M603 8 534 760 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=120980 $D=1
M604 535 759 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=116350 $D=1
M605 536 760 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=120980 $D=1
M606 533 529 535 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=116350 $D=1
M607 534 530 536 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=120980 $D=1
M608 535 106 233 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=116350 $D=1
M609 536 106 234 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=120980 $D=1
M610 237 107 535 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=116350 $D=1
M611 238 107 536 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=120980 $D=1
M612 537 107 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=116350 $D=1
M613 538 107 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=120980 $D=1
M614 8 108 539 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=116350 $D=1
M615 8 108 540 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=120980 $D=1
M616 541 109 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=116350 $D=1
M617 542 109 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=120980 $D=1
M618 8 109 233 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=116350 $D=1
M619 8 109 234 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=120980 $D=1
M620 237 108 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=116350 $D=1
M621 238 108 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=120980 $D=1
M622 8 545 543 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=116350 $D=1
M623 8 546 544 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=120980 $D=1
M624 545 110 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=116350 $D=1
M625 546 110 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=120980 $D=1
M626 761 233 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=116350 $D=1
M627 762 234 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=120980 $D=1
M628 547 543 761 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=116350 $D=1
M629 548 544 762 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=120980 $D=1
M630 8 547 549 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=116350 $D=1
M631 8 548 550 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=120980 $D=1
M632 763 549 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=116350 $D=1
M633 764 550 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=120980 $D=1
M634 547 545 763 8 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=116350 $D=1
M635 548 546 764 8 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=120980 $D=1
M636 8 553 551 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=116350 $D=1
M637 8 554 552 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=120980 $D=1
M638 553 110 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=116350 $D=1
M639 554 110 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=120980 $D=1
M640 765 237 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=116350 $D=1
M641 766 238 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=120980 $D=1
M642 555 551 765 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=116350 $D=1
M643 556 552 766 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=120980 $D=1
M644 8 555 111 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=116350 $D=1
M645 8 556 112 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=120980 $D=1
M646 767 111 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=116350 $D=1
M647 768 112 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=120980 $D=1
M648 555 553 767 8 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=116350 $D=1
M649 556 554 768 8 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=120980 $D=1
M650 557 113 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=116350 $D=1
M651 558 113 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=120980 $D=1
M652 559 557 549 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=116350 $D=1
M653 560 558 550 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=120980 $D=1
M654 114 113 559 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=116350 $D=1
M655 115 113 560 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=120980 $D=1
M656 561 116 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=116350 $D=1
M657 562 116 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=120980 $D=1
M658 563 561 111 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=116350 $D=1
M659 564 562 112 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=120980 $D=1
M660 769 116 563 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=116350 $D=1
M661 770 116 564 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=120980 $D=1
M662 8 111 769 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=116350 $D=1
M663 8 112 770 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=120980 $D=1
M664 565 117 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=116350 $D=1
M665 566 117 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=120980 $D=1
M666 567 565 563 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=116350 $D=1
M667 568 566 564 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=120980 $D=1
M668 9 117 567 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=116350 $D=1
M669 10 117 568 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=120980 $D=1
M670 570 569 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=116350 $D=1
M671 571 118 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=120980 $D=1
M672 8 574 572 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=116350 $D=1
M673 8 575 573 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=120980 $D=1
M674 576 559 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=116350 $D=1
M675 577 560 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=120980 $D=1
M676 574 576 569 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=116350 $D=1
M677 575 577 118 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=120980 $D=1
M678 570 559 574 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=116350 $D=1
M679 571 560 575 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=120980 $D=1
M680 578 572 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=116350 $D=1
M681 579 573 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=120980 $D=1
M682 121 578 567 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=116350 $D=1
M683 569 579 568 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=120980 $D=1
M684 559 572 121 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=116350 $D=1
M685 560 573 569 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=120980 $D=1
M686 580 121 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=116350 $D=1
M687 581 569 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=120980 $D=1
M688 582 572 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=116350 $D=1
M689 583 573 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=120980 $D=1
M690 584 582 580 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=116350 $D=1
M691 585 583 581 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=120980 $D=1
M692 567 572 584 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=116350 $D=1
M693 568 573 585 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=120980 $D=1
M694 586 559 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=116350 $D=1
M695 587 560 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=120980 $D=1
M696 8 567 586 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=116350 $D=1
M697 8 568 587 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=120980 $D=1
M698 588 584 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=116350 $D=1
M699 589 585 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=120980 $D=1
M700 789 559 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=116350 $D=1
M701 790 560 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=120980 $D=1
M702 590 567 789 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=116350 $D=1
M703 591 568 790 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=120980 $D=1
M704 791 559 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=116350 $D=1
M705 792 560 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=120980 $D=1
M706 592 567 791 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=116350 $D=1
M707 593 568 792 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=120980 $D=1
M708 596 559 594 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=116350 $D=1
M709 597 560 595 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=120980 $D=1
M710 594 567 596 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=116350 $D=1
M711 595 568 597 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=120980 $D=1
M712 8 592 594 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=116350 $D=1
M713 8 593 595 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=120980 $D=1
M714 598 124 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=116350 $D=1
M715 599 124 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=120980 $D=1
M716 600 598 586 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=116350 $D=1
M717 601 599 587 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=120980 $D=1
M718 590 124 600 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=116350 $D=1
M719 591 124 601 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=120980 $D=1
M720 602 598 588 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=116350 $D=1
M721 603 599 589 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=120980 $D=1
M722 596 124 602 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=116350 $D=1
M723 597 124 603 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=120980 $D=1
M724 604 125 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=116350 $D=1
M725 605 125 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=120980 $D=1
M726 606 604 602 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=116350 $D=1
M727 607 605 603 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=120980 $D=1
M728 600 125 606 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=116350 $D=1
M729 601 125 607 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=120980 $D=1
M730 11 606 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=116350 $D=1
M731 12 607 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=120980 $D=1
M732 608 126 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=116350 $D=1
M733 609 126 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=120980 $D=1
M734 610 608 127 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=116350 $D=1
M735 611 609 128 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=120980 $D=1
M736 129 126 610 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=116350 $D=1
M737 130 126 611 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=120980 $D=1
M738 612 126 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=116350 $D=1
M739 613 126 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=120980 $D=1
M740 614 612 131 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=116350 $D=1
M741 615 613 132 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=120980 $D=1
M742 133 126 614 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=116350 $D=1
M743 134 126 615 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=120980 $D=1
M744 616 126 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=116350 $D=1
M745 617 126 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=120980 $D=1
M746 618 616 122 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=116350 $D=1
M747 619 617 135 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=120980 $D=1
M748 136 126 618 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=116350 $D=1
M749 137 126 619 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=120980 $D=1
M750 620 126 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=116350 $D=1
M751 621 126 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=120980 $D=1
M752 622 620 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=116350 $D=1
M753 623 621 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=120980 $D=1
M754 138 126 622 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=116350 $D=1
M755 139 126 623 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=120980 $D=1
M756 624 126 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=116350 $D=1
M757 625 126 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=120980 $D=1
M758 626 624 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=116350 $D=1
M759 627 625 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=120980 $D=1
M760 140 126 626 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=116350 $D=1
M761 141 126 627 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=120980 $D=1
M762 8 559 771 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=116350 $D=1
M763 8 560 772 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=120980 $D=1
M764 130 771 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=116350 $D=1
M765 127 772 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=120980 $D=1
M766 628 142 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=116350 $D=1
M767 629 142 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=120980 $D=1
M768 143 628 130 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=116350 $D=1
M769 144 629 127 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=120980 $D=1
M770 610 142 143 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=116350 $D=1
M771 611 142 144 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=120980 $D=1
M772 630 145 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=116350 $D=1
M773 631 145 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=120980 $D=1
M774 146 630 143 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=116350 $D=1
M775 147 631 144 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=120980 $D=1
M776 614 145 146 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=116350 $D=1
M777 615 145 147 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=120980 $D=1
M778 632 148 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=116350 $D=1
M779 633 148 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=120980 $D=1
M780 119 632 146 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=116350 $D=1
M781 120 633 147 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=120980 $D=1
M782 618 148 119 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=116350 $D=1
M783 619 148 120 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=120980 $D=1
M784 634 149 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=116350 $D=1
M785 635 149 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=120980 $D=1
M786 150 634 119 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=116350 $D=1
M787 151 635 120 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=120980 $D=1
M788 622 149 150 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=116350 $D=1
M789 623 149 151 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=120980 $D=1
M790 636 152 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=116350 $D=1
M791 637 152 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=120980 $D=1
M792 209 636 150 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=116350 $D=1
M793 210 637 151 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=120980 $D=1
M794 626 152 209 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=116350 $D=1
M795 627 152 210 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=120980 $D=1
M796 638 153 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=116350 $D=1
M797 639 153 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=120980 $D=1
M798 640 638 111 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=116350 $D=1
M799 641 639 112 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=120980 $D=1
M800 9 153 640 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=116350 $D=1
M801 10 153 641 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=120980 $D=1
M802 793 549 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=116350 $D=1
M803 794 550 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=120980 $D=1
M804 642 640 793 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=116350 $D=1
M805 643 641 794 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=120980 $D=1
M806 646 549 644 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=116350 $D=1
M807 647 550 645 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=120980 $D=1
M808 644 640 646 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=116350 $D=1
M809 645 641 647 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=120980 $D=1
M810 8 642 644 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=116350 $D=1
M811 8 643 645 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=120980 $D=1
M812 795 154 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=116350 $D=1
M813 796 648 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=120980 $D=1
M814 773 646 795 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=116350 $D=1
M815 774 647 796 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=120980 $D=1
M816 648 773 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=116350 $D=1
M817 155 774 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=120980 $D=1
M818 649 549 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=116350 $D=1
M819 650 550 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=120980 $D=1
M820 8 651 649 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=116350 $D=1
M821 8 652 650 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=120980 $D=1
M822 651 640 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=116350 $D=1
M823 652 641 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=120980 $D=1
M824 797 649 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=116350 $D=1
M825 798 650 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=120980 $D=1
M826 653 154 797 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=116350 $D=1
M827 654 648 798 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=120980 $D=1
M828 656 156 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=116350 $D=1
M829 657 655 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=120980 $D=1
M830 799 653 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=116350 $D=1
M831 800 654 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=120980 $D=1
M832 655 656 799 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=116350 $D=1
M833 157 657 800 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=120980 $D=1
M834 659 658 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=116350 $D=1
M835 660 158 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=120980 $D=1
M836 8 663 661 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=116350 $D=1
M837 8 664 662 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=120980 $D=1
M838 665 114 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=116350 $D=1
M839 666 115 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=120980 $D=1
M840 663 665 658 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=116350 $D=1
M841 664 666 158 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=120980 $D=1
M842 659 114 663 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=116350 $D=1
M843 660 115 664 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=120980 $D=1
M844 667 661 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=116350 $D=1
M845 668 662 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=120980 $D=1
M846 159 667 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=116350 $D=1
M847 658 668 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=120980 $D=1
M848 114 661 159 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=116350 $D=1
M849 115 662 658 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=120980 $D=1
M850 669 159 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=116350 $D=1
M851 670 658 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=120980 $D=1
M852 671 661 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=116350 $D=1
M853 672 662 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=120980 $D=1
M854 211 671 669 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=116350 $D=1
M855 212 672 670 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=120980 $D=1
M856 8 661 211 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=116350 $D=1
M857 8 662 212 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=120980 $D=1
M858 673 160 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=116350 $D=1
M859 674 160 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=120980 $D=1
M860 675 673 211 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=116350 $D=1
M861 676 674 212 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=120980 $D=1
M862 11 160 675 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=116350 $D=1
M863 12 160 676 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=120980 $D=1
M864 677 161 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=116350 $D=1
M865 678 161 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=120980 $D=1
M866 679 677 675 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=116350 $D=1
M867 680 678 676 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=120980 $D=1
M868 8 161 679 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=116350 $D=1
M869 8 161 680 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=120980 $D=1
M870 681 110 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=116350 $D=1
M871 682 110 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=120980 $D=1
M872 8 681 683 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=116350 $D=1
M873 8 682 684 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=120980 $D=1
M874 685 110 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=116350 $D=1
M875 686 110 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=120980 $D=1
M876 687 681 679 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=116350 $D=1
M877 688 682 680 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=120980 $D=1
M878 8 687 775 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=116350 $D=1
M879 8 688 776 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=120980 $D=1
M880 689 775 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=116350 $D=1
M881 690 776 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=120980 $D=1
M882 687 683 689 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=116350 $D=1
M883 688 684 690 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=120980 $D=1
M884 691 110 689 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=116350 $D=1
M885 692 110 690 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=120980 $D=1
M886 8 695 693 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=116350 $D=1
M887 8 696 694 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=120980 $D=1
M888 695 110 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=116350 $D=1
M889 696 110 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=120980 $D=1
M890 777 691 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=116350 $D=1
M891 778 692 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=120980 $D=1
M892 697 693 777 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=116350 $D=1
M893 698 694 778 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=120980 $D=1
M894 8 697 114 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=116350 $D=1
M895 8 698 115 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=120980 $D=1
M896 779 114 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=116350 $D=1
M897 780 115 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=120980 $D=1
M898 697 695 779 8 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=116350 $D=1
M899 698 696 780 8 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=120980 $D=1
M900 185 1 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=117600 $D=0
M901 186 1 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=122230 $D=0
M902 187 1 2 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=117600 $D=0
M903 188 1 3 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=122230 $D=0
M904 8 185 187 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=117600 $D=0
M905 8 186 188 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=122230 $D=0
M906 189 1 2 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=117600 $D=0
M907 190 1 3 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=122230 $D=0
M908 2 185 189 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=117600 $D=0
M909 3 186 190 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=122230 $D=0
M910 191 1 2 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=117600 $D=0
M911 192 1 3 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=122230 $D=0
M912 2 185 191 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=117600 $D=0
M913 3 186 192 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=122230 $D=0
M914 195 4 191 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=117600 $D=0
M915 196 4 192 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=122230 $D=0
M916 193 4 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=117600 $D=0
M917 194 4 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=122230 $D=0
M918 197 4 189 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=117600 $D=0
M919 198 4 190 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=122230 $D=0
M920 187 193 197 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=117600 $D=0
M921 188 194 198 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=122230 $D=0
M922 199 5 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=117600 $D=0
M923 200 5 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=122230 $D=0
M924 201 5 197 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=117600 $D=0
M925 202 5 198 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=122230 $D=0
M926 195 199 201 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=117600 $D=0
M927 196 200 202 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=122230 $D=0
M928 203 7 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=117600 $D=0
M929 204 7 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=122230 $D=0
M930 205 7 8 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=117600 $D=0
M931 206 7 8 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=122230 $D=0
M932 9 203 205 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=117600 $D=0
M933 10 204 206 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=122230 $D=0
M934 207 7 11 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=117600 $D=0
M935 208 7 12 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=122230 $D=0
M936 209 203 207 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=117600 $D=0
M937 210 204 208 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=122230 $D=0
M938 213 7 211 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=117600 $D=0
M939 214 7 212 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=122230 $D=0
M940 201 203 213 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=117600 $D=0
M941 202 204 214 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=122230 $D=0
M942 217 13 213 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=117600 $D=0
M943 218 13 214 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=122230 $D=0
M944 215 13 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=117600 $D=0
M945 216 13 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=122230 $D=0
M946 219 13 207 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=117600 $D=0
M947 220 13 208 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=122230 $D=0
M948 205 215 219 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=117600 $D=0
M949 206 216 220 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=122230 $D=0
M950 221 14 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=117600 $D=0
M951 222 14 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=122230 $D=0
M952 223 14 219 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=117600 $D=0
M953 224 14 220 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=122230 $D=0
M954 217 221 223 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=117600 $D=0
M955 218 222 224 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=122230 $D=0
M956 6 15 225 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=117600 $D=0
M957 6 15 226 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=122230 $D=0
M958 227 16 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=117600 $D=0
M959 228 16 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=122230 $D=0
M960 229 225 223 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=117600 $D=0
M961 230 226 224 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=122230 $D=0
M962 6 229 699 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=117600 $D=0
M963 6 230 700 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=122230 $D=0
M964 231 699 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=117600 $D=0
M965 232 700 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=122230 $D=0
M966 229 15 231 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=117600 $D=0
M967 230 15 232 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=122230 $D=0
M968 231 227 233 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=117600 $D=0
M969 232 228 234 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=122230 $D=0
M970 237 235 231 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=117600 $D=0
M971 238 236 232 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=122230 $D=0
M972 235 17 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=117600 $D=0
M973 236 17 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=122230 $D=0
M974 6 18 239 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=117600 $D=0
M975 6 18 240 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=122230 $D=0
M976 241 19 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=117600 $D=0
M977 242 19 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=122230 $D=0
M978 243 239 223 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=117600 $D=0
M979 244 240 224 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=122230 $D=0
M980 6 243 701 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=117600 $D=0
M981 6 244 702 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=122230 $D=0
M982 245 701 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=117600 $D=0
M983 246 702 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=122230 $D=0
M984 243 18 245 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=117600 $D=0
M985 244 18 246 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=122230 $D=0
M986 245 241 233 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=117600 $D=0
M987 246 242 234 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=122230 $D=0
M988 237 247 245 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=117600 $D=0
M989 238 248 246 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=122230 $D=0
M990 247 20 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=117600 $D=0
M991 248 20 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=122230 $D=0
M992 6 21 249 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=117600 $D=0
M993 6 21 250 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=122230 $D=0
M994 251 22 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=117600 $D=0
M995 252 22 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=122230 $D=0
M996 253 249 223 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=117600 $D=0
M997 254 250 224 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=122230 $D=0
M998 6 253 703 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=117600 $D=0
M999 6 254 704 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=122230 $D=0
M1000 255 703 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=117600 $D=0
M1001 256 704 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=122230 $D=0
M1002 253 21 255 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=117600 $D=0
M1003 254 21 256 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=122230 $D=0
M1004 255 251 233 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=117600 $D=0
M1005 256 252 234 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=122230 $D=0
M1006 237 257 255 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=117600 $D=0
M1007 238 258 256 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=122230 $D=0
M1008 257 23 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=117600 $D=0
M1009 258 23 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=122230 $D=0
M1010 6 24 259 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=117600 $D=0
M1011 6 24 260 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=122230 $D=0
M1012 261 25 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=117600 $D=0
M1013 262 25 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=122230 $D=0
M1014 263 259 223 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=117600 $D=0
M1015 264 260 224 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=122230 $D=0
M1016 6 263 705 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=117600 $D=0
M1017 6 264 706 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=122230 $D=0
M1018 265 705 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=117600 $D=0
M1019 266 706 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=122230 $D=0
M1020 263 24 265 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=117600 $D=0
M1021 264 24 266 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=122230 $D=0
M1022 265 261 233 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=117600 $D=0
M1023 266 262 234 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=122230 $D=0
M1024 237 267 265 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=117600 $D=0
M1025 238 268 266 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=122230 $D=0
M1026 267 26 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=117600 $D=0
M1027 268 26 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=122230 $D=0
M1028 6 27 269 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=117600 $D=0
M1029 6 27 270 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=122230 $D=0
M1030 271 28 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=117600 $D=0
M1031 272 28 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=122230 $D=0
M1032 273 269 223 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=117600 $D=0
M1033 274 270 224 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=122230 $D=0
M1034 6 273 707 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=117600 $D=0
M1035 6 274 708 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=122230 $D=0
M1036 275 707 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=117600 $D=0
M1037 276 708 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=122230 $D=0
M1038 273 27 275 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=117600 $D=0
M1039 274 27 276 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=122230 $D=0
M1040 275 271 233 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=117600 $D=0
M1041 276 272 234 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=122230 $D=0
M1042 237 277 275 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=117600 $D=0
M1043 238 278 276 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=122230 $D=0
M1044 277 29 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=117600 $D=0
M1045 278 29 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=122230 $D=0
M1046 6 30 279 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=117600 $D=0
M1047 6 30 280 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=122230 $D=0
M1048 281 31 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=117600 $D=0
M1049 282 31 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=122230 $D=0
M1050 283 279 223 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=117600 $D=0
M1051 284 280 224 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=122230 $D=0
M1052 6 283 709 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=117600 $D=0
M1053 6 284 710 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=122230 $D=0
M1054 285 709 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=117600 $D=0
M1055 286 710 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=122230 $D=0
M1056 283 30 285 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=117600 $D=0
M1057 284 30 286 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=122230 $D=0
M1058 285 281 233 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=117600 $D=0
M1059 286 282 234 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=122230 $D=0
M1060 237 287 285 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=117600 $D=0
M1061 238 288 286 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=122230 $D=0
M1062 287 32 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=117600 $D=0
M1063 288 32 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=122230 $D=0
M1064 6 33 289 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=117600 $D=0
M1065 6 33 290 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=122230 $D=0
M1066 291 34 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=117600 $D=0
M1067 292 34 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=122230 $D=0
M1068 293 289 223 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=117600 $D=0
M1069 294 290 224 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=122230 $D=0
M1070 6 293 711 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=117600 $D=0
M1071 6 294 712 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=122230 $D=0
M1072 295 711 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=117600 $D=0
M1073 296 712 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=122230 $D=0
M1074 293 33 295 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=117600 $D=0
M1075 294 33 296 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=122230 $D=0
M1076 295 291 233 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=117600 $D=0
M1077 296 292 234 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=122230 $D=0
M1078 237 297 295 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=117600 $D=0
M1079 238 298 296 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=122230 $D=0
M1080 297 35 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=117600 $D=0
M1081 298 35 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=122230 $D=0
M1082 6 36 299 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=117600 $D=0
M1083 6 36 300 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=122230 $D=0
M1084 301 37 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=117600 $D=0
M1085 302 37 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=122230 $D=0
M1086 303 299 223 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=117600 $D=0
M1087 304 300 224 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=122230 $D=0
M1088 6 303 713 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=117600 $D=0
M1089 6 304 714 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=122230 $D=0
M1090 305 713 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=117600 $D=0
M1091 306 714 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=122230 $D=0
M1092 303 36 305 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=117600 $D=0
M1093 304 36 306 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=122230 $D=0
M1094 305 301 233 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=117600 $D=0
M1095 306 302 234 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=122230 $D=0
M1096 237 307 305 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=117600 $D=0
M1097 238 308 306 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=122230 $D=0
M1098 307 38 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=117600 $D=0
M1099 308 38 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=122230 $D=0
M1100 6 39 309 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=117600 $D=0
M1101 6 39 310 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=122230 $D=0
M1102 311 40 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=117600 $D=0
M1103 312 40 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=122230 $D=0
M1104 313 309 223 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=117600 $D=0
M1105 314 310 224 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=122230 $D=0
M1106 6 313 715 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=117600 $D=0
M1107 6 314 716 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=122230 $D=0
M1108 315 715 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=117600 $D=0
M1109 316 716 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=122230 $D=0
M1110 313 39 315 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=117600 $D=0
M1111 314 39 316 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=122230 $D=0
M1112 315 311 233 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=117600 $D=0
M1113 316 312 234 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=122230 $D=0
M1114 237 317 315 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=117600 $D=0
M1115 238 318 316 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=122230 $D=0
M1116 317 41 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=117600 $D=0
M1117 318 41 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=122230 $D=0
M1118 6 42 319 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=117600 $D=0
M1119 6 42 320 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=122230 $D=0
M1120 321 43 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=117600 $D=0
M1121 322 43 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=122230 $D=0
M1122 323 319 223 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=117600 $D=0
M1123 324 320 224 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=122230 $D=0
M1124 6 323 717 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=117600 $D=0
M1125 6 324 718 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=122230 $D=0
M1126 325 717 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=117600 $D=0
M1127 326 718 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=122230 $D=0
M1128 323 42 325 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=117600 $D=0
M1129 324 42 326 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=122230 $D=0
M1130 325 321 233 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=117600 $D=0
M1131 326 322 234 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=122230 $D=0
M1132 237 327 325 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=117600 $D=0
M1133 238 328 326 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=122230 $D=0
M1134 327 44 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=117600 $D=0
M1135 328 44 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=122230 $D=0
M1136 6 45 329 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=117600 $D=0
M1137 6 45 330 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=122230 $D=0
M1138 331 46 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=117600 $D=0
M1139 332 46 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=122230 $D=0
M1140 333 329 223 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=117600 $D=0
M1141 334 330 224 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=122230 $D=0
M1142 6 333 719 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=117600 $D=0
M1143 6 334 720 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=122230 $D=0
M1144 335 719 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=117600 $D=0
M1145 336 720 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=122230 $D=0
M1146 333 45 335 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=117600 $D=0
M1147 334 45 336 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=122230 $D=0
M1148 335 331 233 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=117600 $D=0
M1149 336 332 234 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=122230 $D=0
M1150 237 337 335 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=117600 $D=0
M1151 238 338 336 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=122230 $D=0
M1152 337 47 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=117600 $D=0
M1153 338 47 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=122230 $D=0
M1154 6 48 339 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=117600 $D=0
M1155 6 48 340 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=122230 $D=0
M1156 341 49 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=117600 $D=0
M1157 342 49 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=122230 $D=0
M1158 343 339 223 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=117600 $D=0
M1159 344 340 224 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=122230 $D=0
M1160 6 343 721 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=117600 $D=0
M1161 6 344 722 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=122230 $D=0
M1162 345 721 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=117600 $D=0
M1163 346 722 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=122230 $D=0
M1164 343 48 345 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=117600 $D=0
M1165 344 48 346 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=122230 $D=0
M1166 345 341 233 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=117600 $D=0
M1167 346 342 234 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=122230 $D=0
M1168 237 347 345 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=117600 $D=0
M1169 238 348 346 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=122230 $D=0
M1170 347 50 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=117600 $D=0
M1171 348 50 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=122230 $D=0
M1172 6 51 349 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=117600 $D=0
M1173 6 51 350 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=122230 $D=0
M1174 351 52 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=117600 $D=0
M1175 352 52 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=122230 $D=0
M1176 353 349 223 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=117600 $D=0
M1177 354 350 224 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=122230 $D=0
M1178 6 353 723 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=117600 $D=0
M1179 6 354 724 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=122230 $D=0
M1180 355 723 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=117600 $D=0
M1181 356 724 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=122230 $D=0
M1182 353 51 355 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=117600 $D=0
M1183 354 51 356 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=122230 $D=0
M1184 355 351 233 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=117600 $D=0
M1185 356 352 234 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=122230 $D=0
M1186 237 357 355 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=117600 $D=0
M1187 238 358 356 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=122230 $D=0
M1188 357 53 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=117600 $D=0
M1189 358 53 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=122230 $D=0
M1190 6 54 359 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=117600 $D=0
M1191 6 54 360 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=122230 $D=0
M1192 361 55 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=117600 $D=0
M1193 362 55 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=122230 $D=0
M1194 363 359 223 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=117600 $D=0
M1195 364 360 224 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=122230 $D=0
M1196 6 363 725 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=117600 $D=0
M1197 6 364 726 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=122230 $D=0
M1198 365 725 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=117600 $D=0
M1199 366 726 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=122230 $D=0
M1200 363 54 365 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=117600 $D=0
M1201 364 54 366 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=122230 $D=0
M1202 365 361 233 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=117600 $D=0
M1203 366 362 234 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=122230 $D=0
M1204 237 367 365 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=117600 $D=0
M1205 238 368 366 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=122230 $D=0
M1206 367 56 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=117600 $D=0
M1207 368 56 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=122230 $D=0
M1208 6 57 369 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=117600 $D=0
M1209 6 57 370 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=122230 $D=0
M1210 371 58 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=117600 $D=0
M1211 372 58 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=122230 $D=0
M1212 373 369 223 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=117600 $D=0
M1213 374 370 224 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=122230 $D=0
M1214 6 373 727 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=117600 $D=0
M1215 6 374 728 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=122230 $D=0
M1216 375 727 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=117600 $D=0
M1217 376 728 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=122230 $D=0
M1218 373 57 375 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=117600 $D=0
M1219 374 57 376 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=122230 $D=0
M1220 375 371 233 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=117600 $D=0
M1221 376 372 234 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=122230 $D=0
M1222 237 377 375 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=117600 $D=0
M1223 238 378 376 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=122230 $D=0
M1224 377 59 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=117600 $D=0
M1225 378 59 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=122230 $D=0
M1226 6 60 379 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=117600 $D=0
M1227 6 60 380 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=122230 $D=0
M1228 381 61 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=117600 $D=0
M1229 382 61 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=122230 $D=0
M1230 383 379 223 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=117600 $D=0
M1231 384 380 224 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=122230 $D=0
M1232 6 383 729 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=117600 $D=0
M1233 6 384 730 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=122230 $D=0
M1234 385 729 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=117600 $D=0
M1235 386 730 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=122230 $D=0
M1236 383 60 385 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=117600 $D=0
M1237 384 60 386 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=122230 $D=0
M1238 385 381 233 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=117600 $D=0
M1239 386 382 234 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=122230 $D=0
M1240 237 387 385 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=117600 $D=0
M1241 238 388 386 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=122230 $D=0
M1242 387 62 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=117600 $D=0
M1243 388 62 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=122230 $D=0
M1244 6 63 389 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=117600 $D=0
M1245 6 63 390 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=122230 $D=0
M1246 391 64 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=117600 $D=0
M1247 392 64 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=122230 $D=0
M1248 393 389 223 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=117600 $D=0
M1249 394 390 224 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=122230 $D=0
M1250 6 393 731 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=117600 $D=0
M1251 6 394 732 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=122230 $D=0
M1252 395 731 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=117600 $D=0
M1253 396 732 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=122230 $D=0
M1254 393 63 395 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=117600 $D=0
M1255 394 63 396 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=122230 $D=0
M1256 395 391 233 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=117600 $D=0
M1257 396 392 234 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=122230 $D=0
M1258 237 397 395 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=117600 $D=0
M1259 238 398 396 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=122230 $D=0
M1260 397 65 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=117600 $D=0
M1261 398 65 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=122230 $D=0
M1262 6 66 399 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=117600 $D=0
M1263 6 66 400 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=122230 $D=0
M1264 401 67 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=117600 $D=0
M1265 402 67 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=122230 $D=0
M1266 403 399 223 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=117600 $D=0
M1267 404 400 224 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=122230 $D=0
M1268 6 403 733 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=117600 $D=0
M1269 6 404 734 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=122230 $D=0
M1270 405 733 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=117600 $D=0
M1271 406 734 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=122230 $D=0
M1272 403 66 405 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=117600 $D=0
M1273 404 66 406 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=122230 $D=0
M1274 405 401 233 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=117600 $D=0
M1275 406 402 234 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=122230 $D=0
M1276 237 407 405 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=117600 $D=0
M1277 238 408 406 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=122230 $D=0
M1278 407 68 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=117600 $D=0
M1279 408 68 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=122230 $D=0
M1280 6 69 409 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=117600 $D=0
M1281 6 69 410 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=122230 $D=0
M1282 411 70 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=117600 $D=0
M1283 412 70 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=122230 $D=0
M1284 413 409 223 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=117600 $D=0
M1285 414 410 224 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=122230 $D=0
M1286 6 413 735 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=117600 $D=0
M1287 6 414 736 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=122230 $D=0
M1288 415 735 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=117600 $D=0
M1289 416 736 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=122230 $D=0
M1290 413 69 415 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=117600 $D=0
M1291 414 69 416 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=122230 $D=0
M1292 415 411 233 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=117600 $D=0
M1293 416 412 234 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=122230 $D=0
M1294 237 417 415 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=117600 $D=0
M1295 238 418 416 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=122230 $D=0
M1296 417 71 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=117600 $D=0
M1297 418 71 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=122230 $D=0
M1298 6 72 419 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=117600 $D=0
M1299 6 72 420 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=122230 $D=0
M1300 421 73 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=117600 $D=0
M1301 422 73 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=122230 $D=0
M1302 423 419 223 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=117600 $D=0
M1303 424 420 224 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=122230 $D=0
M1304 6 423 737 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=117600 $D=0
M1305 6 424 738 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=122230 $D=0
M1306 425 737 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=117600 $D=0
M1307 426 738 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=122230 $D=0
M1308 423 72 425 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=117600 $D=0
M1309 424 72 426 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=122230 $D=0
M1310 425 421 233 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=117600 $D=0
M1311 426 422 234 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=122230 $D=0
M1312 237 427 425 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=117600 $D=0
M1313 238 428 426 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=122230 $D=0
M1314 427 74 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=117600 $D=0
M1315 428 74 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=122230 $D=0
M1316 6 75 429 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=117600 $D=0
M1317 6 75 430 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=122230 $D=0
M1318 431 76 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=117600 $D=0
M1319 432 76 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=122230 $D=0
M1320 433 429 223 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=117600 $D=0
M1321 434 430 224 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=122230 $D=0
M1322 6 433 739 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=117600 $D=0
M1323 6 434 740 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=122230 $D=0
M1324 435 739 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=117600 $D=0
M1325 436 740 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=122230 $D=0
M1326 433 75 435 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=117600 $D=0
M1327 434 75 436 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=122230 $D=0
M1328 435 431 233 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=117600 $D=0
M1329 436 432 234 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=122230 $D=0
M1330 237 437 435 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=117600 $D=0
M1331 238 438 436 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=122230 $D=0
M1332 437 77 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=117600 $D=0
M1333 438 77 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=122230 $D=0
M1334 6 78 439 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=117600 $D=0
M1335 6 78 440 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=122230 $D=0
M1336 441 79 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=117600 $D=0
M1337 442 79 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=122230 $D=0
M1338 443 439 223 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=117600 $D=0
M1339 444 440 224 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=122230 $D=0
M1340 6 443 741 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=117600 $D=0
M1341 6 444 742 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=122230 $D=0
M1342 445 741 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=117600 $D=0
M1343 446 742 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=122230 $D=0
M1344 443 78 445 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=117600 $D=0
M1345 444 78 446 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=122230 $D=0
M1346 445 441 233 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=117600 $D=0
M1347 446 442 234 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=122230 $D=0
M1348 237 447 445 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=117600 $D=0
M1349 238 448 446 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=122230 $D=0
M1350 447 80 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=117600 $D=0
M1351 448 80 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=122230 $D=0
M1352 6 81 449 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=117600 $D=0
M1353 6 81 450 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=122230 $D=0
M1354 451 82 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=117600 $D=0
M1355 452 82 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=122230 $D=0
M1356 453 449 223 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=117600 $D=0
M1357 454 450 224 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=122230 $D=0
M1358 6 453 743 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=117600 $D=0
M1359 6 454 744 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=122230 $D=0
M1360 455 743 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=117600 $D=0
M1361 456 744 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=122230 $D=0
M1362 453 81 455 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=117600 $D=0
M1363 454 81 456 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=122230 $D=0
M1364 455 451 233 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=117600 $D=0
M1365 456 452 234 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=122230 $D=0
M1366 237 457 455 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=117600 $D=0
M1367 238 458 456 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=122230 $D=0
M1368 457 83 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=117600 $D=0
M1369 458 83 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=122230 $D=0
M1370 6 84 459 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=117600 $D=0
M1371 6 84 460 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=122230 $D=0
M1372 461 85 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=117600 $D=0
M1373 462 85 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=122230 $D=0
M1374 463 459 223 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=117600 $D=0
M1375 464 460 224 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=122230 $D=0
M1376 6 463 745 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=117600 $D=0
M1377 6 464 746 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=122230 $D=0
M1378 465 745 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=117600 $D=0
M1379 466 746 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=122230 $D=0
M1380 463 84 465 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=117600 $D=0
M1381 464 84 466 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=122230 $D=0
M1382 465 461 233 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=117600 $D=0
M1383 466 462 234 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=122230 $D=0
M1384 237 467 465 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=117600 $D=0
M1385 238 468 466 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=122230 $D=0
M1386 467 86 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=117600 $D=0
M1387 468 86 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=122230 $D=0
M1388 6 87 469 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=117600 $D=0
M1389 6 87 470 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=122230 $D=0
M1390 471 88 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=117600 $D=0
M1391 472 88 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=122230 $D=0
M1392 473 469 223 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=117600 $D=0
M1393 474 470 224 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=122230 $D=0
M1394 6 473 747 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=117600 $D=0
M1395 6 474 748 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=122230 $D=0
M1396 475 747 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=117600 $D=0
M1397 476 748 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=122230 $D=0
M1398 473 87 475 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=117600 $D=0
M1399 474 87 476 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=122230 $D=0
M1400 475 471 233 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=117600 $D=0
M1401 476 472 234 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=122230 $D=0
M1402 237 477 475 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=117600 $D=0
M1403 238 478 476 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=122230 $D=0
M1404 477 89 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=117600 $D=0
M1405 478 89 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=122230 $D=0
M1406 6 90 479 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=117600 $D=0
M1407 6 90 480 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=122230 $D=0
M1408 481 91 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=117600 $D=0
M1409 482 91 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=122230 $D=0
M1410 483 479 223 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=117600 $D=0
M1411 484 480 224 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=122230 $D=0
M1412 6 483 749 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=117600 $D=0
M1413 6 484 750 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=122230 $D=0
M1414 485 749 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=117600 $D=0
M1415 486 750 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=122230 $D=0
M1416 483 90 485 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=117600 $D=0
M1417 484 90 486 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=122230 $D=0
M1418 485 481 233 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=117600 $D=0
M1419 486 482 234 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=122230 $D=0
M1420 237 487 485 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=117600 $D=0
M1421 238 488 486 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=122230 $D=0
M1422 487 92 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=117600 $D=0
M1423 488 92 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=122230 $D=0
M1424 6 93 489 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=117600 $D=0
M1425 6 93 490 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=122230 $D=0
M1426 491 94 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=117600 $D=0
M1427 492 94 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=122230 $D=0
M1428 493 489 223 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=117600 $D=0
M1429 494 490 224 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=122230 $D=0
M1430 6 493 751 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=117600 $D=0
M1431 6 494 752 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=122230 $D=0
M1432 495 751 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=117600 $D=0
M1433 496 752 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=122230 $D=0
M1434 493 93 495 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=117600 $D=0
M1435 494 93 496 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=122230 $D=0
M1436 495 491 233 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=117600 $D=0
M1437 496 492 234 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=122230 $D=0
M1438 237 497 495 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=117600 $D=0
M1439 238 498 496 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=122230 $D=0
M1440 497 95 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=117600 $D=0
M1441 498 95 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=122230 $D=0
M1442 6 96 499 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=117600 $D=0
M1443 6 96 500 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=122230 $D=0
M1444 501 97 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=117600 $D=0
M1445 502 97 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=122230 $D=0
M1446 503 499 223 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=117600 $D=0
M1447 504 500 224 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=122230 $D=0
M1448 6 503 753 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=117600 $D=0
M1449 6 504 754 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=122230 $D=0
M1450 505 753 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=117600 $D=0
M1451 506 754 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=122230 $D=0
M1452 503 96 505 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=117600 $D=0
M1453 504 96 506 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=122230 $D=0
M1454 505 501 233 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=117600 $D=0
M1455 506 502 234 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=122230 $D=0
M1456 237 507 505 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=117600 $D=0
M1457 238 508 506 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=122230 $D=0
M1458 507 98 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=117600 $D=0
M1459 508 98 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=122230 $D=0
M1460 6 99 509 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=117600 $D=0
M1461 6 99 510 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=122230 $D=0
M1462 511 100 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=117600 $D=0
M1463 512 100 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=122230 $D=0
M1464 513 509 223 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=117600 $D=0
M1465 514 510 224 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=122230 $D=0
M1466 6 513 755 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=117600 $D=0
M1467 6 514 756 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=122230 $D=0
M1468 515 755 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=117600 $D=0
M1469 516 756 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=122230 $D=0
M1470 513 99 515 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=117600 $D=0
M1471 514 99 516 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=122230 $D=0
M1472 515 511 233 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=117600 $D=0
M1473 516 512 234 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=122230 $D=0
M1474 237 517 515 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=117600 $D=0
M1475 238 518 516 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=122230 $D=0
M1476 517 101 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=117600 $D=0
M1477 518 101 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=122230 $D=0
M1478 6 102 519 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=117600 $D=0
M1479 6 102 520 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=122230 $D=0
M1480 521 103 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=117600 $D=0
M1481 522 103 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=122230 $D=0
M1482 523 519 223 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=117600 $D=0
M1483 524 520 224 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=122230 $D=0
M1484 6 523 757 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=117600 $D=0
M1485 6 524 758 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=122230 $D=0
M1486 525 757 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=117600 $D=0
M1487 526 758 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=122230 $D=0
M1488 523 102 525 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=117600 $D=0
M1489 524 102 526 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=122230 $D=0
M1490 525 521 233 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=117600 $D=0
M1491 526 522 234 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=122230 $D=0
M1492 237 527 525 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=117600 $D=0
M1493 238 528 526 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=122230 $D=0
M1494 527 104 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=117600 $D=0
M1495 528 104 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=122230 $D=0
M1496 6 105 529 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=117600 $D=0
M1497 6 105 530 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=122230 $D=0
M1498 531 106 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=117600 $D=0
M1499 532 106 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=122230 $D=0
M1500 533 529 223 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=117600 $D=0
M1501 534 530 224 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=122230 $D=0
M1502 6 533 759 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=117600 $D=0
M1503 6 534 760 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=122230 $D=0
M1504 535 759 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=117600 $D=0
M1505 536 760 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=122230 $D=0
M1506 533 105 535 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=117600 $D=0
M1507 534 105 536 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=122230 $D=0
M1508 535 531 233 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=117600 $D=0
M1509 536 532 234 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=122230 $D=0
M1510 237 537 535 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=117600 $D=0
M1511 238 538 536 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=122230 $D=0
M1512 537 107 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=117600 $D=0
M1513 538 107 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=122230 $D=0
M1514 6 108 539 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=117600 $D=0
M1515 6 108 540 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=122230 $D=0
M1516 541 109 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=117600 $D=0
M1517 542 109 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=122230 $D=0
M1518 8 541 233 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=117600 $D=0
M1519 8 542 234 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=122230 $D=0
M1520 237 539 8 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=117600 $D=0
M1521 238 540 8 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=122230 $D=0
M1522 6 545 543 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=117600 $D=0
M1523 6 546 544 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=122230 $D=0
M1524 545 110 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=117600 $D=0
M1525 546 110 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=122230 $D=0
M1526 761 233 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=117600 $D=0
M1527 762 234 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=122230 $D=0
M1528 547 545 761 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=117600 $D=0
M1529 548 546 762 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=122230 $D=0
M1530 6 547 549 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=117600 $D=0
M1531 6 548 550 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=122230 $D=0
M1532 763 549 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=117600 $D=0
M1533 764 550 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=122230 $D=0
M1534 547 543 763 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=117600 $D=0
M1535 548 544 764 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=122230 $D=0
M1536 6 553 551 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=117600 $D=0
M1537 6 554 552 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=122230 $D=0
M1538 553 110 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=117600 $D=0
M1539 554 110 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=122230 $D=0
M1540 765 237 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=117600 $D=0
M1541 766 238 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=122230 $D=0
M1542 555 553 765 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=117600 $D=0
M1543 556 554 766 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=122230 $D=0
M1544 6 555 111 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=117600 $D=0
M1545 6 556 112 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=122230 $D=0
M1546 767 111 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=117600 $D=0
M1547 768 112 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=122230 $D=0
M1548 555 551 767 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=117600 $D=0
M1549 556 552 768 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=122230 $D=0
M1550 557 113 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=117600 $D=0
M1551 558 113 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=122230 $D=0
M1552 559 113 549 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=117600 $D=0
M1553 560 113 550 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=122230 $D=0
M1554 114 557 559 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=117600 $D=0
M1555 115 558 560 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=122230 $D=0
M1556 561 116 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=117600 $D=0
M1557 562 116 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=122230 $D=0
M1558 563 116 111 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=117600 $D=0
M1559 564 116 112 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=122230 $D=0
M1560 769 561 563 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=117600 $D=0
M1561 770 562 564 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=122230 $D=0
M1562 6 111 769 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=117600 $D=0
M1563 6 112 770 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=122230 $D=0
M1564 565 117 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=117600 $D=0
M1565 566 117 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=122230 $D=0
M1566 567 117 563 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=117600 $D=0
M1567 568 117 564 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=122230 $D=0
M1568 9 565 567 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=117600 $D=0
M1569 10 566 568 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=122230 $D=0
M1570 570 569 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=117600 $D=0
M1571 571 118 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=122230 $D=0
M1572 6 574 572 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=117600 $D=0
M1573 6 575 573 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=122230 $D=0
M1574 576 559 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=117600 $D=0
M1575 577 560 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=122230 $D=0
M1576 574 559 569 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=117600 $D=0
M1577 575 560 118 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=122230 $D=0
M1578 570 576 574 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=117600 $D=0
M1579 571 577 575 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=122230 $D=0
M1580 578 572 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=117600 $D=0
M1581 579 573 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=122230 $D=0
M1582 121 572 567 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=117600 $D=0
M1583 569 573 568 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=122230 $D=0
M1584 559 578 121 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=117600 $D=0
M1585 560 579 569 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=122230 $D=0
M1586 580 121 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=117600 $D=0
M1587 581 569 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=122230 $D=0
M1588 582 572 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=117600 $D=0
M1589 583 573 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=122230 $D=0
M1590 584 572 580 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=117600 $D=0
M1591 585 573 581 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=122230 $D=0
M1592 567 582 584 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=117600 $D=0
M1593 568 583 585 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=122230 $D=0
M1594 781 559 6 6 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=117240 $D=0
M1595 782 560 6 6 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=121870 $D=0
M1596 586 567 781 6 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=117240 $D=0
M1597 587 568 782 6 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=121870 $D=0
M1598 588 584 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=117600 $D=0
M1599 589 585 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=122230 $D=0
M1600 590 559 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=117600 $D=0
M1601 591 560 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=122230 $D=0
M1602 6 567 590 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=117600 $D=0
M1603 6 568 591 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=122230 $D=0
M1604 592 559 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=117600 $D=0
M1605 593 560 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=122230 $D=0
M1606 6 567 592 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=117600 $D=0
M1607 6 568 593 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=122230 $D=0
M1608 783 559 6 6 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=117420 $D=0
M1609 784 560 6 6 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=122050 $D=0
M1610 596 567 783 6 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=117420 $D=0
M1611 597 568 784 6 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=122050 $D=0
M1612 6 592 596 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=117600 $D=0
M1613 6 593 597 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=122230 $D=0
M1614 598 124 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=117600 $D=0
M1615 599 124 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=122230 $D=0
M1616 600 124 586 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=117600 $D=0
M1617 601 124 587 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=122230 $D=0
M1618 590 598 600 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=117600 $D=0
M1619 591 599 601 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=122230 $D=0
M1620 602 124 588 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=117600 $D=0
M1621 603 124 589 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=122230 $D=0
M1622 596 598 602 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=117600 $D=0
M1623 597 599 603 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=122230 $D=0
M1624 604 125 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=117600 $D=0
M1625 605 125 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=122230 $D=0
M1626 606 125 602 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=117600 $D=0
M1627 607 125 603 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=122230 $D=0
M1628 600 604 606 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=117600 $D=0
M1629 601 605 607 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=122230 $D=0
M1630 11 606 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=117600 $D=0
M1631 12 607 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=122230 $D=0
M1632 608 126 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=117600 $D=0
M1633 609 126 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=122230 $D=0
M1634 610 126 127 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=117600 $D=0
M1635 611 126 128 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=122230 $D=0
M1636 129 608 610 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=117600 $D=0
M1637 130 609 611 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=122230 $D=0
M1638 612 126 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=117600 $D=0
M1639 613 126 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=122230 $D=0
M1640 614 126 131 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=117600 $D=0
M1641 615 126 132 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=122230 $D=0
M1642 133 612 614 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=117600 $D=0
M1643 134 613 615 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=122230 $D=0
M1644 616 126 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=117600 $D=0
M1645 617 126 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=122230 $D=0
M1646 618 126 122 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=117600 $D=0
M1647 619 126 135 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=122230 $D=0
M1648 136 616 618 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=117600 $D=0
M1649 137 617 619 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=122230 $D=0
M1650 620 126 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=117600 $D=0
M1651 621 126 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=122230 $D=0
M1652 622 126 8 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=117600 $D=0
M1653 623 126 8 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=122230 $D=0
M1654 138 620 622 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=117600 $D=0
M1655 139 621 623 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=122230 $D=0
M1656 624 126 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=117600 $D=0
M1657 625 126 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=122230 $D=0
M1658 626 126 8 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=117600 $D=0
M1659 627 126 8 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=122230 $D=0
M1660 140 624 626 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=117600 $D=0
M1661 141 625 627 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=122230 $D=0
M1662 6 559 771 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=117600 $D=0
M1663 6 560 772 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=122230 $D=0
M1664 130 771 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=117600 $D=0
M1665 127 772 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=122230 $D=0
M1666 628 142 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=117600 $D=0
M1667 629 142 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=122230 $D=0
M1668 143 142 130 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=117600 $D=0
M1669 144 142 127 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=122230 $D=0
M1670 610 628 143 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=117600 $D=0
M1671 611 629 144 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=122230 $D=0
M1672 630 145 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=117600 $D=0
M1673 631 145 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=122230 $D=0
M1674 146 145 143 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=117600 $D=0
M1675 147 145 144 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=122230 $D=0
M1676 614 630 146 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=117600 $D=0
M1677 615 631 147 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=122230 $D=0
M1678 632 148 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=117600 $D=0
M1679 633 148 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=122230 $D=0
M1680 119 148 146 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=117600 $D=0
M1681 120 148 147 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=122230 $D=0
M1682 618 632 119 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=117600 $D=0
M1683 619 633 120 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=122230 $D=0
M1684 634 149 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=117600 $D=0
M1685 635 149 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=122230 $D=0
M1686 150 149 119 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=117600 $D=0
M1687 151 149 120 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=122230 $D=0
M1688 622 634 150 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=117600 $D=0
M1689 623 635 151 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=122230 $D=0
M1690 636 152 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=117600 $D=0
M1691 637 152 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=122230 $D=0
M1692 209 152 150 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=117600 $D=0
M1693 210 152 151 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=122230 $D=0
M1694 626 636 209 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=117600 $D=0
M1695 627 637 210 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=122230 $D=0
M1696 638 153 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=117600 $D=0
M1697 639 153 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=122230 $D=0
M1698 640 153 111 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=117600 $D=0
M1699 641 153 112 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=122230 $D=0
M1700 9 638 640 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=117600 $D=0
M1701 10 639 641 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=122230 $D=0
M1702 642 549 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=117600 $D=0
M1703 643 550 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=122230 $D=0
M1704 6 640 642 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=117600 $D=0
M1705 6 641 643 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=122230 $D=0
M1706 785 549 6 6 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=117420 $D=0
M1707 786 550 6 6 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=122050 $D=0
M1708 646 640 785 6 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=117420 $D=0
M1709 647 641 786 6 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=122050 $D=0
M1710 6 642 646 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=117600 $D=0
M1711 6 643 647 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=122230 $D=0
M1712 773 154 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=117600 $D=0
M1713 774 648 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=122230 $D=0
M1714 6 646 773 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=117600 $D=0
M1715 6 647 774 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=122230 $D=0
M1716 648 773 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=117600 $D=0
M1717 155 774 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=122230 $D=0
M1718 787 549 6 6 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=117240 $D=0
M1719 788 550 6 6 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=121870 $D=0
M1720 649 651 787 6 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=117240 $D=0
M1721 650 652 788 6 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=121870 $D=0
M1722 651 640 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=117600 $D=0
M1723 652 641 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=122230 $D=0
M1724 653 649 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=117600 $D=0
M1725 654 650 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=122230 $D=0
M1726 6 154 653 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=117600 $D=0
M1727 6 648 654 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=122230 $D=0
M1728 656 156 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=117600 $D=0
M1729 657 655 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=122230 $D=0
M1730 655 653 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=117600 $D=0
M1731 157 654 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=122230 $D=0
M1732 6 656 655 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=117600 $D=0
M1733 6 657 157 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=122230 $D=0
M1734 659 658 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=117600 $D=0
M1735 660 158 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=122230 $D=0
M1736 6 663 661 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=117600 $D=0
M1737 6 664 662 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=122230 $D=0
M1738 665 114 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=117600 $D=0
M1739 666 115 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=122230 $D=0
M1740 663 114 658 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=117600 $D=0
M1741 664 115 158 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=122230 $D=0
M1742 659 665 663 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=117600 $D=0
M1743 660 666 664 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=122230 $D=0
M1744 667 661 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=117600 $D=0
M1745 668 662 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=122230 $D=0
M1746 159 661 8 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=117600 $D=0
M1747 658 662 8 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=122230 $D=0
M1748 114 667 159 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=117600 $D=0
M1749 115 668 658 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=122230 $D=0
M1750 669 159 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=117600 $D=0
M1751 670 658 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=122230 $D=0
M1752 671 661 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=117600 $D=0
M1753 672 662 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=122230 $D=0
M1754 211 661 669 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=117600 $D=0
M1755 212 662 670 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=122230 $D=0
M1756 8 671 211 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=117600 $D=0
M1757 8 672 212 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=122230 $D=0
M1758 673 160 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=117600 $D=0
M1759 674 160 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=122230 $D=0
M1760 675 160 211 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=117600 $D=0
M1761 676 160 212 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=122230 $D=0
M1762 11 673 675 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=117600 $D=0
M1763 12 674 676 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=122230 $D=0
M1764 677 161 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=117600 $D=0
M1765 678 161 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=122230 $D=0
M1766 679 161 675 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=117600 $D=0
M1767 680 161 676 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=122230 $D=0
M1768 8 677 679 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=117600 $D=0
M1769 8 678 680 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=122230 $D=0
M1770 681 110 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=117600 $D=0
M1771 682 110 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=122230 $D=0
M1772 6 681 683 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=117600 $D=0
M1773 6 682 684 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=122230 $D=0
M1774 685 110 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=117600 $D=0
M1775 686 110 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=122230 $D=0
M1776 687 683 679 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=117600 $D=0
M1777 688 684 680 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=122230 $D=0
M1778 6 687 775 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=117600 $D=0
M1779 6 688 776 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=122230 $D=0
M1780 689 775 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=117600 $D=0
M1781 690 776 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=122230 $D=0
M1782 687 681 689 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=117600 $D=0
M1783 688 682 690 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=122230 $D=0
M1784 691 685 689 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=117600 $D=0
M1785 692 686 690 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=122230 $D=0
M1786 6 695 693 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=117600 $D=0
M1787 6 696 694 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=122230 $D=0
M1788 695 110 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=117600 $D=0
M1789 696 110 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=122230 $D=0
M1790 777 691 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=117600 $D=0
M1791 778 692 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=122230 $D=0
M1792 697 695 777 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=117600 $D=0
M1793 698 696 778 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=122230 $D=0
M1794 6 697 114 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=117600 $D=0
M1795 6 698 115 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=122230 $D=0
M1796 779 114 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=117600 $D=0
M1797 780 115 6 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=122230 $D=0
M1798 697 693 779 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=117600 $D=0
M1799 698 694 780 6 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=122230 $D=0
.ENDS
***************************************
.SUBCKT ICV_27 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161
** N=807 EP=161 IP=1514 FDC=1800
M0 192 1 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=107090 $D=1
M1 193 1 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=111720 $D=1
M2 194 192 2 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=107090 $D=1
M3 195 193 3 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=111720 $D=1
M4 4 1 194 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=107090 $D=1
M5 4 1 195 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=111720 $D=1
M6 196 192 3 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=107090 $D=1
M7 197 193 3 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=111720 $D=1
M8 2 1 196 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=107090 $D=1
M9 3 1 197 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=111720 $D=1
M10 198 192 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=107090 $D=1
M11 199 193 3 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=111720 $D=1
M12 2 1 198 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=107090 $D=1
M13 3 1 199 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=111720 $D=1
M14 202 200 198 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=107090 $D=1
M15 203 201 199 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=111720 $D=1
M16 200 5 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=107090 $D=1
M17 201 5 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=111720 $D=1
M18 204 200 196 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=107090 $D=1
M19 205 201 197 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=111720 $D=1
M20 194 5 204 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=107090 $D=1
M21 195 5 205 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=111720 $D=1
M22 206 6 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=107090 $D=1
M23 207 6 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=111720 $D=1
M24 208 206 204 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=107090 $D=1
M25 209 207 205 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=111720 $D=1
M26 202 6 208 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=107090 $D=1
M27 203 6 209 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=111720 $D=1
M28 210 8 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=107090 $D=1
M29 211 8 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=111720 $D=1
M30 212 210 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=107090 $D=1
M31 213 211 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=111720 $D=1
M32 9 8 212 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=107090 $D=1
M33 10 8 213 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=111720 $D=1
M34 214 210 11 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=107090 $D=1
M35 215 211 12 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=111720 $D=1
M36 216 8 214 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=107090 $D=1
M37 217 8 215 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=111720 $D=1
M38 220 210 218 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=107090 $D=1
M39 221 211 219 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=111720 $D=1
M40 208 8 220 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=107090 $D=1
M41 209 8 221 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=111720 $D=1
M42 224 222 220 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=107090 $D=1
M43 225 223 221 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=111720 $D=1
M44 222 13 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=107090 $D=1
M45 223 13 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=111720 $D=1
M46 226 222 214 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=107090 $D=1
M47 227 223 215 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=111720 $D=1
M48 212 13 226 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=107090 $D=1
M49 213 13 227 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=111720 $D=1
M50 228 14 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=107090 $D=1
M51 229 14 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=111720 $D=1
M52 230 228 226 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=107090 $D=1
M53 231 229 227 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=111720 $D=1
M54 224 14 230 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=107090 $D=1
M55 225 14 231 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=111720 $D=1
M56 4 15 232 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=107090 $D=1
M57 4 15 233 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=111720 $D=1
M58 234 16 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=107090 $D=1
M59 235 16 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=111720 $D=1
M60 236 15 230 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=107090 $D=1
M61 237 15 231 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=111720 $D=1
M62 4 236 706 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=107090 $D=1
M63 4 237 707 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=111720 $D=1
M64 238 706 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=107090 $D=1
M65 239 707 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=111720 $D=1
M66 236 232 238 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=107090 $D=1
M67 237 233 239 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=111720 $D=1
M68 238 16 240 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=107090 $D=1
M69 239 16 241 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=111720 $D=1
M70 244 17 238 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=107090 $D=1
M71 245 17 239 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=111720 $D=1
M72 242 17 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=107090 $D=1
M73 243 17 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=111720 $D=1
M74 4 18 246 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=107090 $D=1
M75 4 18 247 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=111720 $D=1
M76 248 19 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=107090 $D=1
M77 249 19 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=111720 $D=1
M78 250 18 230 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=107090 $D=1
M79 251 18 231 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=111720 $D=1
M80 4 250 708 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=107090 $D=1
M81 4 251 709 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=111720 $D=1
M82 252 708 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=107090 $D=1
M83 253 709 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=111720 $D=1
M84 250 246 252 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=107090 $D=1
M85 251 247 253 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=111720 $D=1
M86 252 19 240 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=107090 $D=1
M87 253 19 241 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=111720 $D=1
M88 244 20 252 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=107090 $D=1
M89 245 20 253 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=111720 $D=1
M90 254 20 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=107090 $D=1
M91 255 20 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=111720 $D=1
M92 4 21 256 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=107090 $D=1
M93 4 21 257 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=111720 $D=1
M94 258 22 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=107090 $D=1
M95 259 22 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=111720 $D=1
M96 260 21 230 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=107090 $D=1
M97 261 21 231 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=111720 $D=1
M98 4 260 710 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=107090 $D=1
M99 4 261 711 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=111720 $D=1
M100 262 710 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=107090 $D=1
M101 263 711 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=111720 $D=1
M102 260 256 262 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=107090 $D=1
M103 261 257 263 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=111720 $D=1
M104 262 22 240 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=107090 $D=1
M105 263 22 241 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=111720 $D=1
M106 244 23 262 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=107090 $D=1
M107 245 23 263 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=111720 $D=1
M108 264 23 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=107090 $D=1
M109 265 23 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=111720 $D=1
M110 4 24 266 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=107090 $D=1
M111 4 24 267 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=111720 $D=1
M112 268 25 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=107090 $D=1
M113 269 25 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=111720 $D=1
M114 270 24 230 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=107090 $D=1
M115 271 24 231 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=111720 $D=1
M116 4 270 712 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=107090 $D=1
M117 4 271 713 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=111720 $D=1
M118 272 712 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=107090 $D=1
M119 273 713 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=111720 $D=1
M120 270 266 272 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=107090 $D=1
M121 271 267 273 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=111720 $D=1
M122 272 25 240 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=107090 $D=1
M123 273 25 241 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=111720 $D=1
M124 244 26 272 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=107090 $D=1
M125 245 26 273 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=111720 $D=1
M126 274 26 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=107090 $D=1
M127 275 26 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=111720 $D=1
M128 4 27 276 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=107090 $D=1
M129 4 27 277 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=111720 $D=1
M130 278 28 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=107090 $D=1
M131 279 28 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=111720 $D=1
M132 280 27 230 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=107090 $D=1
M133 281 27 231 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=111720 $D=1
M134 4 280 714 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=107090 $D=1
M135 4 281 715 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=111720 $D=1
M136 282 714 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=107090 $D=1
M137 283 715 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=111720 $D=1
M138 280 276 282 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=107090 $D=1
M139 281 277 283 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=111720 $D=1
M140 282 28 240 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=107090 $D=1
M141 283 28 241 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=111720 $D=1
M142 244 29 282 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=107090 $D=1
M143 245 29 283 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=111720 $D=1
M144 284 29 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=107090 $D=1
M145 285 29 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=111720 $D=1
M146 4 30 286 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=107090 $D=1
M147 4 30 287 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=111720 $D=1
M148 288 31 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=107090 $D=1
M149 289 31 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=111720 $D=1
M150 290 30 230 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=107090 $D=1
M151 291 30 231 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=111720 $D=1
M152 4 290 716 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=107090 $D=1
M153 4 291 717 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=111720 $D=1
M154 292 716 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=107090 $D=1
M155 293 717 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=111720 $D=1
M156 290 286 292 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=107090 $D=1
M157 291 287 293 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=111720 $D=1
M158 292 31 240 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=107090 $D=1
M159 293 31 241 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=111720 $D=1
M160 244 32 292 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=107090 $D=1
M161 245 32 293 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=111720 $D=1
M162 294 32 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=107090 $D=1
M163 295 32 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=111720 $D=1
M164 4 33 296 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=107090 $D=1
M165 4 33 297 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=111720 $D=1
M166 298 34 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=107090 $D=1
M167 299 34 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=111720 $D=1
M168 300 33 230 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=107090 $D=1
M169 301 33 231 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=111720 $D=1
M170 4 300 718 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=107090 $D=1
M171 4 301 719 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=111720 $D=1
M172 302 718 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=107090 $D=1
M173 303 719 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=111720 $D=1
M174 300 296 302 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=107090 $D=1
M175 301 297 303 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=111720 $D=1
M176 302 34 240 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=107090 $D=1
M177 303 34 241 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=111720 $D=1
M178 244 35 302 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=107090 $D=1
M179 245 35 303 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=111720 $D=1
M180 304 35 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=107090 $D=1
M181 305 35 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=111720 $D=1
M182 4 36 306 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=107090 $D=1
M183 4 36 307 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=111720 $D=1
M184 308 37 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=107090 $D=1
M185 309 37 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=111720 $D=1
M186 310 36 230 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=107090 $D=1
M187 311 36 231 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=111720 $D=1
M188 4 310 720 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=107090 $D=1
M189 4 311 721 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=111720 $D=1
M190 312 720 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=107090 $D=1
M191 313 721 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=111720 $D=1
M192 310 306 312 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=107090 $D=1
M193 311 307 313 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=111720 $D=1
M194 312 37 240 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=107090 $D=1
M195 313 37 241 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=111720 $D=1
M196 244 38 312 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=107090 $D=1
M197 245 38 313 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=111720 $D=1
M198 314 38 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=107090 $D=1
M199 315 38 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=111720 $D=1
M200 4 39 316 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=107090 $D=1
M201 4 39 317 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=111720 $D=1
M202 318 40 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=107090 $D=1
M203 319 40 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=111720 $D=1
M204 320 39 230 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=107090 $D=1
M205 321 39 231 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=111720 $D=1
M206 4 320 722 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=107090 $D=1
M207 4 321 723 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=111720 $D=1
M208 322 722 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=107090 $D=1
M209 323 723 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=111720 $D=1
M210 320 316 322 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=107090 $D=1
M211 321 317 323 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=111720 $D=1
M212 322 40 240 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=107090 $D=1
M213 323 40 241 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=111720 $D=1
M214 244 41 322 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=107090 $D=1
M215 245 41 323 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=111720 $D=1
M216 324 41 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=107090 $D=1
M217 325 41 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=111720 $D=1
M218 4 42 326 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=107090 $D=1
M219 4 42 327 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=111720 $D=1
M220 328 43 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=107090 $D=1
M221 329 43 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=111720 $D=1
M222 330 42 230 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=107090 $D=1
M223 331 42 231 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=111720 $D=1
M224 4 330 724 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=107090 $D=1
M225 4 331 725 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=111720 $D=1
M226 332 724 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=107090 $D=1
M227 333 725 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=111720 $D=1
M228 330 326 332 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=107090 $D=1
M229 331 327 333 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=111720 $D=1
M230 332 43 240 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=107090 $D=1
M231 333 43 241 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=111720 $D=1
M232 244 44 332 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=107090 $D=1
M233 245 44 333 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=111720 $D=1
M234 334 44 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=107090 $D=1
M235 335 44 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=111720 $D=1
M236 4 45 336 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=107090 $D=1
M237 4 45 337 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=111720 $D=1
M238 338 46 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=107090 $D=1
M239 339 46 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=111720 $D=1
M240 340 45 230 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=107090 $D=1
M241 341 45 231 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=111720 $D=1
M242 4 340 726 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=107090 $D=1
M243 4 341 727 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=111720 $D=1
M244 342 726 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=107090 $D=1
M245 343 727 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=111720 $D=1
M246 340 336 342 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=107090 $D=1
M247 341 337 343 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=111720 $D=1
M248 342 46 240 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=107090 $D=1
M249 343 46 241 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=111720 $D=1
M250 244 47 342 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=107090 $D=1
M251 245 47 343 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=111720 $D=1
M252 344 47 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=107090 $D=1
M253 345 47 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=111720 $D=1
M254 4 48 346 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=107090 $D=1
M255 4 48 347 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=111720 $D=1
M256 348 49 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=107090 $D=1
M257 349 49 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=111720 $D=1
M258 350 48 230 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=107090 $D=1
M259 351 48 231 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=111720 $D=1
M260 4 350 728 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=107090 $D=1
M261 4 351 729 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=111720 $D=1
M262 352 728 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=107090 $D=1
M263 353 729 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=111720 $D=1
M264 350 346 352 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=107090 $D=1
M265 351 347 353 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=111720 $D=1
M266 352 49 240 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=107090 $D=1
M267 353 49 241 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=111720 $D=1
M268 244 50 352 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=107090 $D=1
M269 245 50 353 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=111720 $D=1
M270 354 50 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=107090 $D=1
M271 355 50 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=111720 $D=1
M272 4 51 356 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=107090 $D=1
M273 4 51 357 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=111720 $D=1
M274 358 52 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=107090 $D=1
M275 359 52 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=111720 $D=1
M276 360 51 230 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=107090 $D=1
M277 361 51 231 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=111720 $D=1
M278 4 360 730 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=107090 $D=1
M279 4 361 731 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=111720 $D=1
M280 362 730 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=107090 $D=1
M281 363 731 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=111720 $D=1
M282 360 356 362 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=107090 $D=1
M283 361 357 363 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=111720 $D=1
M284 362 52 240 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=107090 $D=1
M285 363 52 241 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=111720 $D=1
M286 244 53 362 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=107090 $D=1
M287 245 53 363 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=111720 $D=1
M288 364 53 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=107090 $D=1
M289 365 53 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=111720 $D=1
M290 4 54 366 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=107090 $D=1
M291 4 54 367 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=111720 $D=1
M292 368 55 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=107090 $D=1
M293 369 55 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=111720 $D=1
M294 370 54 230 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=107090 $D=1
M295 371 54 231 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=111720 $D=1
M296 4 370 732 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=107090 $D=1
M297 4 371 733 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=111720 $D=1
M298 372 732 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=107090 $D=1
M299 373 733 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=111720 $D=1
M300 370 366 372 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=107090 $D=1
M301 371 367 373 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=111720 $D=1
M302 372 55 240 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=107090 $D=1
M303 373 55 241 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=111720 $D=1
M304 244 56 372 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=107090 $D=1
M305 245 56 373 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=111720 $D=1
M306 374 56 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=107090 $D=1
M307 375 56 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=111720 $D=1
M308 4 57 376 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=107090 $D=1
M309 4 57 377 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=111720 $D=1
M310 378 58 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=107090 $D=1
M311 379 58 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=111720 $D=1
M312 380 57 230 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=107090 $D=1
M313 381 57 231 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=111720 $D=1
M314 4 380 734 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=107090 $D=1
M315 4 381 735 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=111720 $D=1
M316 382 734 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=107090 $D=1
M317 383 735 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=111720 $D=1
M318 380 376 382 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=107090 $D=1
M319 381 377 383 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=111720 $D=1
M320 382 58 240 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=107090 $D=1
M321 383 58 241 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=111720 $D=1
M322 244 59 382 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=107090 $D=1
M323 245 59 383 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=111720 $D=1
M324 384 59 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=107090 $D=1
M325 385 59 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=111720 $D=1
M326 4 60 386 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=107090 $D=1
M327 4 60 387 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=111720 $D=1
M328 388 61 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=107090 $D=1
M329 389 61 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=111720 $D=1
M330 390 60 230 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=107090 $D=1
M331 391 60 231 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=111720 $D=1
M332 4 390 736 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=107090 $D=1
M333 4 391 737 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=111720 $D=1
M334 392 736 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=107090 $D=1
M335 393 737 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=111720 $D=1
M336 390 386 392 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=107090 $D=1
M337 391 387 393 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=111720 $D=1
M338 392 61 240 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=107090 $D=1
M339 393 61 241 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=111720 $D=1
M340 244 62 392 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=107090 $D=1
M341 245 62 393 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=111720 $D=1
M342 394 62 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=107090 $D=1
M343 395 62 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=111720 $D=1
M344 4 63 396 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=107090 $D=1
M345 4 63 397 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=111720 $D=1
M346 398 64 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=107090 $D=1
M347 399 64 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=111720 $D=1
M348 400 63 230 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=107090 $D=1
M349 401 63 231 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=111720 $D=1
M350 4 400 738 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=107090 $D=1
M351 4 401 739 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=111720 $D=1
M352 402 738 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=107090 $D=1
M353 403 739 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=111720 $D=1
M354 400 396 402 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=107090 $D=1
M355 401 397 403 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=111720 $D=1
M356 402 64 240 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=107090 $D=1
M357 403 64 241 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=111720 $D=1
M358 244 65 402 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=107090 $D=1
M359 245 65 403 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=111720 $D=1
M360 404 65 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=107090 $D=1
M361 405 65 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=111720 $D=1
M362 4 66 406 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=107090 $D=1
M363 4 66 407 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=111720 $D=1
M364 408 67 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=107090 $D=1
M365 409 67 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=111720 $D=1
M366 410 66 230 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=107090 $D=1
M367 411 66 231 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=111720 $D=1
M368 4 410 740 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=107090 $D=1
M369 4 411 741 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=111720 $D=1
M370 412 740 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=107090 $D=1
M371 413 741 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=111720 $D=1
M372 410 406 412 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=107090 $D=1
M373 411 407 413 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=111720 $D=1
M374 412 67 240 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=107090 $D=1
M375 413 67 241 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=111720 $D=1
M376 244 68 412 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=107090 $D=1
M377 245 68 413 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=111720 $D=1
M378 414 68 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=107090 $D=1
M379 415 68 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=111720 $D=1
M380 4 69 416 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=107090 $D=1
M381 4 69 417 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=111720 $D=1
M382 418 70 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=107090 $D=1
M383 419 70 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=111720 $D=1
M384 420 69 230 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=107090 $D=1
M385 421 69 231 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=111720 $D=1
M386 4 420 742 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=107090 $D=1
M387 4 421 743 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=111720 $D=1
M388 422 742 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=107090 $D=1
M389 423 743 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=111720 $D=1
M390 420 416 422 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=107090 $D=1
M391 421 417 423 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=111720 $D=1
M392 422 70 240 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=107090 $D=1
M393 423 70 241 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=111720 $D=1
M394 244 71 422 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=107090 $D=1
M395 245 71 423 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=111720 $D=1
M396 424 71 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=107090 $D=1
M397 425 71 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=111720 $D=1
M398 4 72 426 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=107090 $D=1
M399 4 72 427 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=111720 $D=1
M400 428 73 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=107090 $D=1
M401 429 73 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=111720 $D=1
M402 430 72 230 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=107090 $D=1
M403 431 72 231 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=111720 $D=1
M404 4 430 744 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=107090 $D=1
M405 4 431 745 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=111720 $D=1
M406 432 744 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=107090 $D=1
M407 433 745 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=111720 $D=1
M408 430 426 432 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=107090 $D=1
M409 431 427 433 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=111720 $D=1
M410 432 73 240 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=107090 $D=1
M411 433 73 241 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=111720 $D=1
M412 244 74 432 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=107090 $D=1
M413 245 74 433 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=111720 $D=1
M414 434 74 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=107090 $D=1
M415 435 74 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=111720 $D=1
M416 4 75 436 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=107090 $D=1
M417 4 75 437 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=111720 $D=1
M418 438 76 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=107090 $D=1
M419 439 76 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=111720 $D=1
M420 440 75 230 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=107090 $D=1
M421 441 75 231 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=111720 $D=1
M422 4 440 746 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=107090 $D=1
M423 4 441 747 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=111720 $D=1
M424 442 746 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=107090 $D=1
M425 443 747 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=111720 $D=1
M426 440 436 442 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=107090 $D=1
M427 441 437 443 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=111720 $D=1
M428 442 76 240 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=107090 $D=1
M429 443 76 241 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=111720 $D=1
M430 244 77 442 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=107090 $D=1
M431 245 77 443 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=111720 $D=1
M432 444 77 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=107090 $D=1
M433 445 77 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=111720 $D=1
M434 4 78 446 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=107090 $D=1
M435 4 78 447 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=111720 $D=1
M436 448 79 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=107090 $D=1
M437 449 79 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=111720 $D=1
M438 450 78 230 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=107090 $D=1
M439 451 78 231 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=111720 $D=1
M440 4 450 748 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=107090 $D=1
M441 4 451 749 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=111720 $D=1
M442 452 748 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=107090 $D=1
M443 453 749 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=111720 $D=1
M444 450 446 452 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=107090 $D=1
M445 451 447 453 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=111720 $D=1
M446 452 79 240 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=107090 $D=1
M447 453 79 241 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=111720 $D=1
M448 244 80 452 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=107090 $D=1
M449 245 80 453 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=111720 $D=1
M450 454 80 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=107090 $D=1
M451 455 80 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=111720 $D=1
M452 4 81 456 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=107090 $D=1
M453 4 81 457 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=111720 $D=1
M454 458 82 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=107090 $D=1
M455 459 82 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=111720 $D=1
M456 460 81 230 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=107090 $D=1
M457 461 81 231 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=111720 $D=1
M458 4 460 750 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=107090 $D=1
M459 4 461 751 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=111720 $D=1
M460 462 750 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=107090 $D=1
M461 463 751 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=111720 $D=1
M462 460 456 462 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=107090 $D=1
M463 461 457 463 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=111720 $D=1
M464 462 82 240 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=107090 $D=1
M465 463 82 241 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=111720 $D=1
M466 244 83 462 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=107090 $D=1
M467 245 83 463 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=111720 $D=1
M468 464 83 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=107090 $D=1
M469 465 83 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=111720 $D=1
M470 4 84 466 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=107090 $D=1
M471 4 84 467 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=111720 $D=1
M472 468 85 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=107090 $D=1
M473 469 85 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=111720 $D=1
M474 470 84 230 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=107090 $D=1
M475 471 84 231 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=111720 $D=1
M476 4 470 752 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=107090 $D=1
M477 4 471 753 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=111720 $D=1
M478 472 752 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=107090 $D=1
M479 473 753 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=111720 $D=1
M480 470 466 472 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=107090 $D=1
M481 471 467 473 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=111720 $D=1
M482 472 85 240 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=107090 $D=1
M483 473 85 241 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=111720 $D=1
M484 244 86 472 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=107090 $D=1
M485 245 86 473 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=111720 $D=1
M486 474 86 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=107090 $D=1
M487 475 86 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=111720 $D=1
M488 4 87 476 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=107090 $D=1
M489 4 87 477 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=111720 $D=1
M490 478 88 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=107090 $D=1
M491 479 88 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=111720 $D=1
M492 480 87 230 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=107090 $D=1
M493 481 87 231 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=111720 $D=1
M494 4 480 754 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=107090 $D=1
M495 4 481 755 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=111720 $D=1
M496 482 754 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=107090 $D=1
M497 483 755 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=111720 $D=1
M498 480 476 482 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=107090 $D=1
M499 481 477 483 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=111720 $D=1
M500 482 88 240 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=107090 $D=1
M501 483 88 241 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=111720 $D=1
M502 244 89 482 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=107090 $D=1
M503 245 89 483 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=111720 $D=1
M504 484 89 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=107090 $D=1
M505 485 89 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=111720 $D=1
M506 4 90 486 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=107090 $D=1
M507 4 90 487 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=111720 $D=1
M508 488 91 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=107090 $D=1
M509 489 91 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=111720 $D=1
M510 490 90 230 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=107090 $D=1
M511 491 90 231 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=111720 $D=1
M512 4 490 756 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=107090 $D=1
M513 4 491 757 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=111720 $D=1
M514 492 756 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=107090 $D=1
M515 493 757 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=111720 $D=1
M516 490 486 492 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=107090 $D=1
M517 491 487 493 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=111720 $D=1
M518 492 91 240 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=107090 $D=1
M519 493 91 241 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=111720 $D=1
M520 244 92 492 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=107090 $D=1
M521 245 92 493 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=111720 $D=1
M522 494 92 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=107090 $D=1
M523 495 92 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=111720 $D=1
M524 4 93 496 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=107090 $D=1
M525 4 93 497 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=111720 $D=1
M526 498 94 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=107090 $D=1
M527 499 94 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=111720 $D=1
M528 500 93 230 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=107090 $D=1
M529 501 93 231 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=111720 $D=1
M530 4 500 758 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=107090 $D=1
M531 4 501 759 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=111720 $D=1
M532 502 758 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=107090 $D=1
M533 503 759 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=111720 $D=1
M534 500 496 502 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=107090 $D=1
M535 501 497 503 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=111720 $D=1
M536 502 94 240 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=107090 $D=1
M537 503 94 241 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=111720 $D=1
M538 244 95 502 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=107090 $D=1
M539 245 95 503 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=111720 $D=1
M540 504 95 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=107090 $D=1
M541 505 95 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=111720 $D=1
M542 4 96 506 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=107090 $D=1
M543 4 96 507 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=111720 $D=1
M544 508 97 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=107090 $D=1
M545 509 97 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=111720 $D=1
M546 510 96 230 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=107090 $D=1
M547 511 96 231 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=111720 $D=1
M548 4 510 760 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=107090 $D=1
M549 4 511 761 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=111720 $D=1
M550 512 760 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=107090 $D=1
M551 513 761 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=111720 $D=1
M552 510 506 512 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=107090 $D=1
M553 511 507 513 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=111720 $D=1
M554 512 97 240 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=107090 $D=1
M555 513 97 241 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=111720 $D=1
M556 244 98 512 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=107090 $D=1
M557 245 98 513 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=111720 $D=1
M558 514 98 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=107090 $D=1
M559 515 98 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=111720 $D=1
M560 4 99 516 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=107090 $D=1
M561 4 99 517 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=111720 $D=1
M562 518 100 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=107090 $D=1
M563 519 100 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=111720 $D=1
M564 520 99 230 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=107090 $D=1
M565 521 99 231 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=111720 $D=1
M566 4 520 762 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=107090 $D=1
M567 4 521 763 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=111720 $D=1
M568 522 762 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=107090 $D=1
M569 523 763 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=111720 $D=1
M570 520 516 522 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=107090 $D=1
M571 521 517 523 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=111720 $D=1
M572 522 100 240 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=107090 $D=1
M573 523 100 241 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=111720 $D=1
M574 244 101 522 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=107090 $D=1
M575 245 101 523 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=111720 $D=1
M576 524 101 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=107090 $D=1
M577 525 101 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=111720 $D=1
M578 4 102 526 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=107090 $D=1
M579 4 102 527 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=111720 $D=1
M580 528 103 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=107090 $D=1
M581 529 103 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=111720 $D=1
M582 530 102 230 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=107090 $D=1
M583 531 102 231 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=111720 $D=1
M584 4 530 764 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=107090 $D=1
M585 4 531 765 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=111720 $D=1
M586 532 764 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=107090 $D=1
M587 533 765 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=111720 $D=1
M588 530 526 532 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=107090 $D=1
M589 531 527 533 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=111720 $D=1
M590 532 103 240 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=107090 $D=1
M591 533 103 241 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=111720 $D=1
M592 244 104 532 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=107090 $D=1
M593 245 104 533 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=111720 $D=1
M594 534 104 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=107090 $D=1
M595 535 104 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=111720 $D=1
M596 4 105 536 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=107090 $D=1
M597 4 105 537 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=111720 $D=1
M598 538 106 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=107090 $D=1
M599 539 106 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=111720 $D=1
M600 540 105 230 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=107090 $D=1
M601 541 105 231 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=111720 $D=1
M602 4 540 766 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=107090 $D=1
M603 4 541 767 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=111720 $D=1
M604 542 766 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=107090 $D=1
M605 543 767 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=111720 $D=1
M606 540 536 542 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=107090 $D=1
M607 541 537 543 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=111720 $D=1
M608 542 106 240 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=107090 $D=1
M609 543 106 241 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=111720 $D=1
M610 244 107 542 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=107090 $D=1
M611 245 107 543 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=111720 $D=1
M612 544 107 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=107090 $D=1
M613 545 107 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=111720 $D=1
M614 4 108 546 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=107090 $D=1
M615 4 108 547 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=111720 $D=1
M616 548 109 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=107090 $D=1
M617 549 109 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=111720 $D=1
M618 4 109 240 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=107090 $D=1
M619 4 109 241 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=111720 $D=1
M620 244 108 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=107090 $D=1
M621 245 108 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=111720 $D=1
M622 4 552 550 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=107090 $D=1
M623 4 553 551 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=111720 $D=1
M624 552 110 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=107090 $D=1
M625 553 110 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=111720 $D=1
M626 768 240 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=107090 $D=1
M627 769 241 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=111720 $D=1
M628 554 550 768 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=107090 $D=1
M629 555 551 769 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=111720 $D=1
M630 4 554 556 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=107090 $D=1
M631 4 555 557 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=111720 $D=1
M632 770 556 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=107090 $D=1
M633 771 557 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=111720 $D=1
M634 554 552 770 4 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=107090 $D=1
M635 555 553 771 4 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=111720 $D=1
M636 4 560 558 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=107090 $D=1
M637 4 561 559 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=111720 $D=1
M638 560 110 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=107090 $D=1
M639 561 110 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=111720 $D=1
M640 772 244 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=107090 $D=1
M641 773 245 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=111720 $D=1
M642 562 558 772 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=107090 $D=1
M643 563 559 773 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=111720 $D=1
M644 4 562 111 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=107090 $D=1
M645 4 563 112 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=111720 $D=1
M646 774 111 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=107090 $D=1
M647 775 112 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=111720 $D=1
M648 562 560 774 4 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=107090 $D=1
M649 563 561 775 4 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=111720 $D=1
M650 564 113 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=107090 $D=1
M651 565 113 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=111720 $D=1
M652 566 564 556 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=107090 $D=1
M653 567 565 557 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=111720 $D=1
M654 114 113 566 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=107090 $D=1
M655 115 113 567 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=111720 $D=1
M656 568 116 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=107090 $D=1
M657 569 116 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=111720 $D=1
M658 570 568 111 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=107090 $D=1
M659 571 569 112 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=111720 $D=1
M660 776 116 570 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=107090 $D=1
M661 777 116 571 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=111720 $D=1
M662 4 111 776 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=107090 $D=1
M663 4 112 777 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=111720 $D=1
M664 572 118 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=107090 $D=1
M665 573 118 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=111720 $D=1
M666 574 572 570 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=107090 $D=1
M667 575 573 571 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=111720 $D=1
M668 9 118 574 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=107090 $D=1
M669 10 118 575 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=111720 $D=1
M670 577 576 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=107090 $D=1
M671 578 120 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=111720 $D=1
M672 4 581 579 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=107090 $D=1
M673 4 582 580 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=111720 $D=1
M674 583 566 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=107090 $D=1
M675 584 567 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=111720 $D=1
M676 581 583 576 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=107090 $D=1
M677 582 584 120 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=111720 $D=1
M678 577 566 581 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=107090 $D=1
M679 578 567 582 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=111720 $D=1
M680 585 579 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=107090 $D=1
M681 586 580 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=111720 $D=1
M682 124 585 574 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=107090 $D=1
M683 576 586 575 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=111720 $D=1
M684 566 579 124 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=107090 $D=1
M685 567 580 576 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=111720 $D=1
M686 587 124 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=107090 $D=1
M687 588 576 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=111720 $D=1
M688 589 579 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=107090 $D=1
M689 590 580 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=111720 $D=1
M690 591 589 587 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=107090 $D=1
M691 592 590 588 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=111720 $D=1
M692 574 579 591 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=107090 $D=1
M693 575 580 592 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=111720 $D=1
M694 593 566 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=107090 $D=1
M695 594 567 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=111720 $D=1
M696 4 574 593 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=107090 $D=1
M697 4 575 594 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=111720 $D=1
M698 595 591 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=107090 $D=1
M699 596 592 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=111720 $D=1
M700 796 566 4 4 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=107090 $D=1
M701 797 567 4 4 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=111720 $D=1
M702 597 574 796 4 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=107090 $D=1
M703 598 575 797 4 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=111720 $D=1
M704 798 566 4 4 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=107090 $D=1
M705 799 567 4 4 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=111720 $D=1
M706 599 574 798 4 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=107090 $D=1
M707 600 575 799 4 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=111720 $D=1
M708 603 566 601 4 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=107090 $D=1
M709 604 567 602 4 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=111720 $D=1
M710 601 574 603 4 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=107090 $D=1
M711 602 575 604 4 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=111720 $D=1
M712 4 599 601 4 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=107090 $D=1
M713 4 600 602 4 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=111720 $D=1
M714 605 126 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=107090 $D=1
M715 606 126 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=111720 $D=1
M716 607 605 593 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=107090 $D=1
M717 608 606 594 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=111720 $D=1
M718 597 126 607 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=107090 $D=1
M719 598 126 608 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=111720 $D=1
M720 609 605 595 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=107090 $D=1
M721 610 606 596 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=111720 $D=1
M722 603 126 609 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=107090 $D=1
M723 604 126 610 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=111720 $D=1
M724 611 127 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=107090 $D=1
M725 612 127 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=111720 $D=1
M726 613 611 609 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=107090 $D=1
M727 614 612 610 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=111720 $D=1
M728 607 127 613 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=107090 $D=1
M729 608 127 614 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=111720 $D=1
M730 11 613 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=107090 $D=1
M731 12 614 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=111720 $D=1
M732 615 128 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=107090 $D=1
M733 616 128 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=111720 $D=1
M734 617 615 129 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=107090 $D=1
M735 618 616 130 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=111720 $D=1
M736 131 128 617 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=107090 $D=1
M737 132 128 618 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=111720 $D=1
M738 619 128 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=107090 $D=1
M739 620 128 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=111720 $D=1
M740 621 619 133 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=107090 $D=1
M741 622 620 134 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=111720 $D=1
M742 135 128 621 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=107090 $D=1
M743 136 128 622 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=111720 $D=1
M744 623 128 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=107090 $D=1
M745 624 128 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=111720 $D=1
M746 625 623 137 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=107090 $D=1
M747 626 624 138 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=111720 $D=1
M748 117 128 625 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=107090 $D=1
M749 123 128 626 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=111720 $D=1
M750 627 128 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=107090 $D=1
M751 628 128 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=111720 $D=1
M752 629 627 139 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=107090 $D=1
M753 630 628 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=111720 $D=1
M754 119 128 629 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=107090 $D=1
M755 140 128 630 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=111720 $D=1
M756 631 128 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=107090 $D=1
M757 632 128 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=111720 $D=1
M758 633 631 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=107090 $D=1
M759 634 632 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=111720 $D=1
M760 141 128 633 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=107090 $D=1
M761 142 128 634 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=111720 $D=1
M762 4 566 778 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=107090 $D=1
M763 4 567 779 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=111720 $D=1
M764 132 778 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=107090 $D=1
M765 129 779 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=111720 $D=1
M766 635 143 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=107090 $D=1
M767 636 143 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=111720 $D=1
M768 144 635 132 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=107090 $D=1
M769 145 636 129 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=111720 $D=1
M770 617 143 144 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=107090 $D=1
M771 618 143 145 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=111720 $D=1
M772 637 146 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=107090 $D=1
M773 638 146 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=111720 $D=1
M774 125 637 144 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=107090 $D=1
M775 147 638 145 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=111720 $D=1
M776 621 146 125 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=107090 $D=1
M777 622 146 147 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=111720 $D=1
M778 639 148 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=107090 $D=1
M779 640 148 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=111720 $D=1
M780 121 639 125 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=107090 $D=1
M781 122 640 147 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=111720 $D=1
M782 625 148 121 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=107090 $D=1
M783 626 148 122 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=111720 $D=1
M784 641 149 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=107090 $D=1
M785 642 149 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=111720 $D=1
M786 150 641 121 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=107090 $D=1
M787 151 642 122 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=111720 $D=1
M788 629 149 150 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=107090 $D=1
M789 630 149 151 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=111720 $D=1
M790 643 152 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=107090 $D=1
M791 644 152 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=111720 $D=1
M792 216 643 150 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=107090 $D=1
M793 217 644 151 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=111720 $D=1
M794 633 152 216 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=107090 $D=1
M795 634 152 217 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=111720 $D=1
M796 645 153 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=107090 $D=1
M797 646 153 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=111720 $D=1
M798 647 645 111 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=107090 $D=1
M799 648 646 112 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=111720 $D=1
M800 9 153 647 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=107090 $D=1
M801 10 153 648 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=111720 $D=1
M802 800 556 4 4 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=107090 $D=1
M803 801 557 4 4 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=111720 $D=1
M804 649 647 800 4 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=107090 $D=1
M805 650 648 801 4 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=111720 $D=1
M806 653 556 651 4 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=107090 $D=1
M807 654 557 652 4 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=111720 $D=1
M808 651 647 653 4 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=107090 $D=1
M809 652 648 654 4 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=111720 $D=1
M810 4 649 651 4 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=107090 $D=1
M811 4 650 652 4 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=111720 $D=1
M812 802 154 4 4 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=107090 $D=1
M813 803 655 4 4 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=111720 $D=1
M814 780 653 802 4 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=107090 $D=1
M815 781 654 803 4 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=111720 $D=1
M816 655 780 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=107090 $D=1
M817 155 781 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=111720 $D=1
M818 656 556 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=107090 $D=1
M819 657 557 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=111720 $D=1
M820 4 658 656 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=107090 $D=1
M821 4 659 657 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=111720 $D=1
M822 658 647 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=107090 $D=1
M823 659 648 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=111720 $D=1
M824 804 656 4 4 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=107090 $D=1
M825 805 657 4 4 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=111720 $D=1
M826 660 154 804 4 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=107090 $D=1
M827 661 655 805 4 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=111720 $D=1
M828 663 156 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=107090 $D=1
M829 664 662 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=111720 $D=1
M830 806 660 4 4 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=107090 $D=1
M831 807 661 4 4 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=111720 $D=1
M832 662 663 806 4 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=107090 $D=1
M833 157 664 807 4 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=111720 $D=1
M834 666 665 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=107090 $D=1
M835 667 158 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=111720 $D=1
M836 4 670 668 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=107090 $D=1
M837 4 671 669 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=111720 $D=1
M838 672 114 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=107090 $D=1
M839 673 115 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=111720 $D=1
M840 670 672 665 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=107090 $D=1
M841 671 673 158 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=111720 $D=1
M842 666 114 670 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=107090 $D=1
M843 667 115 671 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=111720 $D=1
M844 674 668 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=107090 $D=1
M845 675 669 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=111720 $D=1
M846 159 674 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=107090 $D=1
M847 665 675 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=111720 $D=1
M848 114 668 159 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=107090 $D=1
M849 115 669 665 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=111720 $D=1
M850 676 159 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=107090 $D=1
M851 677 665 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=111720 $D=1
M852 678 668 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=107090 $D=1
M853 679 669 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=111720 $D=1
M854 218 678 676 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=107090 $D=1
M855 219 679 677 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=111720 $D=1
M856 4 668 218 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=107090 $D=1
M857 4 669 219 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=111720 $D=1
M858 680 160 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=107090 $D=1
M859 681 160 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=111720 $D=1
M860 682 680 218 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=107090 $D=1
M861 683 681 219 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=111720 $D=1
M862 11 160 682 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=107090 $D=1
M863 12 160 683 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=111720 $D=1
M864 684 161 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=107090 $D=1
M865 685 161 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=111720 $D=1
M866 686 684 682 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=107090 $D=1
M867 687 685 683 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=111720 $D=1
M868 4 161 686 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=107090 $D=1
M869 4 161 687 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=111720 $D=1
M870 688 110 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=107090 $D=1
M871 689 110 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=111720 $D=1
M872 4 688 690 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=107090 $D=1
M873 4 689 691 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=111720 $D=1
M874 692 110 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=107090 $D=1
M875 693 110 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=111720 $D=1
M876 694 688 686 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=107090 $D=1
M877 695 689 687 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=111720 $D=1
M878 4 694 782 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=107090 $D=1
M879 4 695 783 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=111720 $D=1
M880 696 782 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=107090 $D=1
M881 697 783 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=111720 $D=1
M882 694 690 696 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=107090 $D=1
M883 695 691 697 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=111720 $D=1
M884 698 110 696 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=107090 $D=1
M885 699 110 697 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=111720 $D=1
M886 4 702 700 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=107090 $D=1
M887 4 703 701 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=111720 $D=1
M888 702 110 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=107090 $D=1
M889 703 110 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=111720 $D=1
M890 784 698 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=107090 $D=1
M891 785 699 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=111720 $D=1
M892 704 700 784 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=107090 $D=1
M893 705 701 785 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=111720 $D=1
M894 4 704 114 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=107090 $D=1
M895 4 705 115 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=111720 $D=1
M896 786 114 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=107090 $D=1
M897 787 115 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=111720 $D=1
M898 704 702 786 4 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=107090 $D=1
M899 705 703 787 4 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=111720 $D=1
M900 192 1 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=108340 $D=0
M901 193 1 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=112970 $D=0
M902 194 1 2 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=108340 $D=0
M903 195 1 3 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=112970 $D=0
M904 4 192 194 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=108340 $D=0
M905 4 193 195 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=112970 $D=0
M906 196 1 3 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=108340 $D=0
M907 197 1 3 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=112970 $D=0
M908 2 192 196 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=108340 $D=0
M909 3 193 197 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=112970 $D=0
M910 198 1 4 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=108340 $D=0
M911 199 1 3 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=112970 $D=0
M912 2 192 198 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=108340 $D=0
M913 3 193 199 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=112970 $D=0
M914 202 5 198 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=108340 $D=0
M915 203 5 199 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=112970 $D=0
M916 200 5 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=108340 $D=0
M917 201 5 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=112970 $D=0
M918 204 5 196 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=108340 $D=0
M919 205 5 197 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=112970 $D=0
M920 194 200 204 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=108340 $D=0
M921 195 201 205 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=112970 $D=0
M922 206 6 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=108340 $D=0
M923 207 6 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=112970 $D=0
M924 208 6 204 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=108340 $D=0
M925 209 6 205 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=112970 $D=0
M926 202 206 208 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=108340 $D=0
M927 203 207 209 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=112970 $D=0
M928 210 8 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=108340 $D=0
M929 211 8 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=112970 $D=0
M930 212 8 4 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=108340 $D=0
M931 213 8 4 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=112970 $D=0
M932 9 210 212 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=108340 $D=0
M933 10 211 213 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=112970 $D=0
M934 214 8 11 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=108340 $D=0
M935 215 8 12 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=112970 $D=0
M936 216 210 214 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=108340 $D=0
M937 217 211 215 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=112970 $D=0
M938 220 8 218 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=108340 $D=0
M939 221 8 219 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=112970 $D=0
M940 208 210 220 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=108340 $D=0
M941 209 211 221 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=112970 $D=0
M942 224 13 220 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=108340 $D=0
M943 225 13 221 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=112970 $D=0
M944 222 13 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=108340 $D=0
M945 223 13 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=112970 $D=0
M946 226 13 214 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=108340 $D=0
M947 227 13 215 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=112970 $D=0
M948 212 222 226 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=108340 $D=0
M949 213 223 227 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=112970 $D=0
M950 228 14 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=108340 $D=0
M951 229 14 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=112970 $D=0
M952 230 14 226 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=108340 $D=0
M953 231 14 227 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=112970 $D=0
M954 224 228 230 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=108340 $D=0
M955 225 229 231 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=112970 $D=0
M956 7 15 232 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=108340 $D=0
M957 7 15 233 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=112970 $D=0
M958 234 16 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=108340 $D=0
M959 235 16 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=112970 $D=0
M960 236 232 230 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=108340 $D=0
M961 237 233 231 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=112970 $D=0
M962 7 236 706 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=108340 $D=0
M963 7 237 707 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=112970 $D=0
M964 238 706 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=108340 $D=0
M965 239 707 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=112970 $D=0
M966 236 15 238 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=108340 $D=0
M967 237 15 239 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=112970 $D=0
M968 238 234 240 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=108340 $D=0
M969 239 235 241 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=112970 $D=0
M970 244 242 238 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=108340 $D=0
M971 245 243 239 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=112970 $D=0
M972 242 17 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=108340 $D=0
M973 243 17 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=112970 $D=0
M974 7 18 246 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=108340 $D=0
M975 7 18 247 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=112970 $D=0
M976 248 19 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=108340 $D=0
M977 249 19 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=112970 $D=0
M978 250 246 230 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=108340 $D=0
M979 251 247 231 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=112970 $D=0
M980 7 250 708 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=108340 $D=0
M981 7 251 709 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=112970 $D=0
M982 252 708 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=108340 $D=0
M983 253 709 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=112970 $D=0
M984 250 18 252 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=108340 $D=0
M985 251 18 253 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=112970 $D=0
M986 252 248 240 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=108340 $D=0
M987 253 249 241 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=112970 $D=0
M988 244 254 252 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=108340 $D=0
M989 245 255 253 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=112970 $D=0
M990 254 20 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=108340 $D=0
M991 255 20 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=112970 $D=0
M992 7 21 256 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=108340 $D=0
M993 7 21 257 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=112970 $D=0
M994 258 22 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=108340 $D=0
M995 259 22 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=112970 $D=0
M996 260 256 230 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=108340 $D=0
M997 261 257 231 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=112970 $D=0
M998 7 260 710 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=108340 $D=0
M999 7 261 711 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=112970 $D=0
M1000 262 710 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=108340 $D=0
M1001 263 711 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=112970 $D=0
M1002 260 21 262 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=108340 $D=0
M1003 261 21 263 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=112970 $D=0
M1004 262 258 240 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=108340 $D=0
M1005 263 259 241 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=112970 $D=0
M1006 244 264 262 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=108340 $D=0
M1007 245 265 263 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=112970 $D=0
M1008 264 23 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=108340 $D=0
M1009 265 23 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=112970 $D=0
M1010 7 24 266 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=108340 $D=0
M1011 7 24 267 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=112970 $D=0
M1012 268 25 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=108340 $D=0
M1013 269 25 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=112970 $D=0
M1014 270 266 230 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=108340 $D=0
M1015 271 267 231 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=112970 $D=0
M1016 7 270 712 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=108340 $D=0
M1017 7 271 713 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=112970 $D=0
M1018 272 712 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=108340 $D=0
M1019 273 713 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=112970 $D=0
M1020 270 24 272 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=108340 $D=0
M1021 271 24 273 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=112970 $D=0
M1022 272 268 240 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=108340 $D=0
M1023 273 269 241 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=112970 $D=0
M1024 244 274 272 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=108340 $D=0
M1025 245 275 273 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=112970 $D=0
M1026 274 26 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=108340 $D=0
M1027 275 26 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=112970 $D=0
M1028 7 27 276 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=108340 $D=0
M1029 7 27 277 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=112970 $D=0
M1030 278 28 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=108340 $D=0
M1031 279 28 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=112970 $D=0
M1032 280 276 230 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=108340 $D=0
M1033 281 277 231 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=112970 $D=0
M1034 7 280 714 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=108340 $D=0
M1035 7 281 715 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=112970 $D=0
M1036 282 714 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=108340 $D=0
M1037 283 715 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=112970 $D=0
M1038 280 27 282 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=108340 $D=0
M1039 281 27 283 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=112970 $D=0
M1040 282 278 240 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=108340 $D=0
M1041 283 279 241 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=112970 $D=0
M1042 244 284 282 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=108340 $D=0
M1043 245 285 283 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=112970 $D=0
M1044 284 29 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=108340 $D=0
M1045 285 29 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=112970 $D=0
M1046 7 30 286 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=108340 $D=0
M1047 7 30 287 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=112970 $D=0
M1048 288 31 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=108340 $D=0
M1049 289 31 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=112970 $D=0
M1050 290 286 230 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=108340 $D=0
M1051 291 287 231 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=112970 $D=0
M1052 7 290 716 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=108340 $D=0
M1053 7 291 717 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=112970 $D=0
M1054 292 716 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=108340 $D=0
M1055 293 717 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=112970 $D=0
M1056 290 30 292 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=108340 $D=0
M1057 291 30 293 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=112970 $D=0
M1058 292 288 240 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=108340 $D=0
M1059 293 289 241 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=112970 $D=0
M1060 244 294 292 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=108340 $D=0
M1061 245 295 293 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=112970 $D=0
M1062 294 32 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=108340 $D=0
M1063 295 32 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=112970 $D=0
M1064 7 33 296 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=108340 $D=0
M1065 7 33 297 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=112970 $D=0
M1066 298 34 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=108340 $D=0
M1067 299 34 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=112970 $D=0
M1068 300 296 230 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=108340 $D=0
M1069 301 297 231 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=112970 $D=0
M1070 7 300 718 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=108340 $D=0
M1071 7 301 719 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=112970 $D=0
M1072 302 718 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=108340 $D=0
M1073 303 719 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=112970 $D=0
M1074 300 33 302 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=108340 $D=0
M1075 301 33 303 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=112970 $D=0
M1076 302 298 240 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=108340 $D=0
M1077 303 299 241 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=112970 $D=0
M1078 244 304 302 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=108340 $D=0
M1079 245 305 303 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=112970 $D=0
M1080 304 35 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=108340 $D=0
M1081 305 35 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=112970 $D=0
M1082 7 36 306 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=108340 $D=0
M1083 7 36 307 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=112970 $D=0
M1084 308 37 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=108340 $D=0
M1085 309 37 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=112970 $D=0
M1086 310 306 230 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=108340 $D=0
M1087 311 307 231 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=112970 $D=0
M1088 7 310 720 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=108340 $D=0
M1089 7 311 721 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=112970 $D=0
M1090 312 720 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=108340 $D=0
M1091 313 721 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=112970 $D=0
M1092 310 36 312 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=108340 $D=0
M1093 311 36 313 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=112970 $D=0
M1094 312 308 240 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=108340 $D=0
M1095 313 309 241 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=112970 $D=0
M1096 244 314 312 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=108340 $D=0
M1097 245 315 313 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=112970 $D=0
M1098 314 38 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=108340 $D=0
M1099 315 38 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=112970 $D=0
M1100 7 39 316 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=108340 $D=0
M1101 7 39 317 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=112970 $D=0
M1102 318 40 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=108340 $D=0
M1103 319 40 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=112970 $D=0
M1104 320 316 230 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=108340 $D=0
M1105 321 317 231 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=112970 $D=0
M1106 7 320 722 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=108340 $D=0
M1107 7 321 723 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=112970 $D=0
M1108 322 722 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=108340 $D=0
M1109 323 723 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=112970 $D=0
M1110 320 39 322 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=108340 $D=0
M1111 321 39 323 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=112970 $D=0
M1112 322 318 240 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=108340 $D=0
M1113 323 319 241 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=112970 $D=0
M1114 244 324 322 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=108340 $D=0
M1115 245 325 323 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=112970 $D=0
M1116 324 41 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=108340 $D=0
M1117 325 41 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=112970 $D=0
M1118 7 42 326 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=108340 $D=0
M1119 7 42 327 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=112970 $D=0
M1120 328 43 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=108340 $D=0
M1121 329 43 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=112970 $D=0
M1122 330 326 230 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=108340 $D=0
M1123 331 327 231 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=112970 $D=0
M1124 7 330 724 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=108340 $D=0
M1125 7 331 725 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=112970 $D=0
M1126 332 724 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=108340 $D=0
M1127 333 725 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=112970 $D=0
M1128 330 42 332 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=108340 $D=0
M1129 331 42 333 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=112970 $D=0
M1130 332 328 240 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=108340 $D=0
M1131 333 329 241 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=112970 $D=0
M1132 244 334 332 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=108340 $D=0
M1133 245 335 333 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=112970 $D=0
M1134 334 44 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=108340 $D=0
M1135 335 44 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=112970 $D=0
M1136 7 45 336 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=108340 $D=0
M1137 7 45 337 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=112970 $D=0
M1138 338 46 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=108340 $D=0
M1139 339 46 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=112970 $D=0
M1140 340 336 230 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=108340 $D=0
M1141 341 337 231 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=112970 $D=0
M1142 7 340 726 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=108340 $D=0
M1143 7 341 727 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=112970 $D=0
M1144 342 726 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=108340 $D=0
M1145 343 727 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=112970 $D=0
M1146 340 45 342 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=108340 $D=0
M1147 341 45 343 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=112970 $D=0
M1148 342 338 240 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=108340 $D=0
M1149 343 339 241 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=112970 $D=0
M1150 244 344 342 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=108340 $D=0
M1151 245 345 343 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=112970 $D=0
M1152 344 47 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=108340 $D=0
M1153 345 47 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=112970 $D=0
M1154 7 48 346 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=108340 $D=0
M1155 7 48 347 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=112970 $D=0
M1156 348 49 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=108340 $D=0
M1157 349 49 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=112970 $D=0
M1158 350 346 230 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=108340 $D=0
M1159 351 347 231 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=112970 $D=0
M1160 7 350 728 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=108340 $D=0
M1161 7 351 729 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=112970 $D=0
M1162 352 728 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=108340 $D=0
M1163 353 729 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=112970 $D=0
M1164 350 48 352 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=108340 $D=0
M1165 351 48 353 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=112970 $D=0
M1166 352 348 240 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=108340 $D=0
M1167 353 349 241 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=112970 $D=0
M1168 244 354 352 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=108340 $D=0
M1169 245 355 353 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=112970 $D=0
M1170 354 50 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=108340 $D=0
M1171 355 50 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=112970 $D=0
M1172 7 51 356 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=108340 $D=0
M1173 7 51 357 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=112970 $D=0
M1174 358 52 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=108340 $D=0
M1175 359 52 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=112970 $D=0
M1176 360 356 230 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=108340 $D=0
M1177 361 357 231 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=112970 $D=0
M1178 7 360 730 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=108340 $D=0
M1179 7 361 731 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=112970 $D=0
M1180 362 730 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=108340 $D=0
M1181 363 731 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=112970 $D=0
M1182 360 51 362 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=108340 $D=0
M1183 361 51 363 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=112970 $D=0
M1184 362 358 240 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=108340 $D=0
M1185 363 359 241 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=112970 $D=0
M1186 244 364 362 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=108340 $D=0
M1187 245 365 363 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=112970 $D=0
M1188 364 53 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=108340 $D=0
M1189 365 53 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=112970 $D=0
M1190 7 54 366 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=108340 $D=0
M1191 7 54 367 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=112970 $D=0
M1192 368 55 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=108340 $D=0
M1193 369 55 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=112970 $D=0
M1194 370 366 230 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=108340 $D=0
M1195 371 367 231 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=112970 $D=0
M1196 7 370 732 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=108340 $D=0
M1197 7 371 733 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=112970 $D=0
M1198 372 732 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=108340 $D=0
M1199 373 733 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=112970 $D=0
M1200 370 54 372 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=108340 $D=0
M1201 371 54 373 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=112970 $D=0
M1202 372 368 240 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=108340 $D=0
M1203 373 369 241 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=112970 $D=0
M1204 244 374 372 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=108340 $D=0
M1205 245 375 373 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=112970 $D=0
M1206 374 56 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=108340 $D=0
M1207 375 56 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=112970 $D=0
M1208 7 57 376 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=108340 $D=0
M1209 7 57 377 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=112970 $D=0
M1210 378 58 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=108340 $D=0
M1211 379 58 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=112970 $D=0
M1212 380 376 230 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=108340 $D=0
M1213 381 377 231 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=112970 $D=0
M1214 7 380 734 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=108340 $D=0
M1215 7 381 735 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=112970 $D=0
M1216 382 734 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=108340 $D=0
M1217 383 735 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=112970 $D=0
M1218 380 57 382 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=108340 $D=0
M1219 381 57 383 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=112970 $D=0
M1220 382 378 240 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=108340 $D=0
M1221 383 379 241 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=112970 $D=0
M1222 244 384 382 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=108340 $D=0
M1223 245 385 383 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=112970 $D=0
M1224 384 59 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=108340 $D=0
M1225 385 59 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=112970 $D=0
M1226 7 60 386 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=108340 $D=0
M1227 7 60 387 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=112970 $D=0
M1228 388 61 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=108340 $D=0
M1229 389 61 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=112970 $D=0
M1230 390 386 230 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=108340 $D=0
M1231 391 387 231 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=112970 $D=0
M1232 7 390 736 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=108340 $D=0
M1233 7 391 737 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=112970 $D=0
M1234 392 736 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=108340 $D=0
M1235 393 737 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=112970 $D=0
M1236 390 60 392 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=108340 $D=0
M1237 391 60 393 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=112970 $D=0
M1238 392 388 240 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=108340 $D=0
M1239 393 389 241 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=112970 $D=0
M1240 244 394 392 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=108340 $D=0
M1241 245 395 393 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=112970 $D=0
M1242 394 62 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=108340 $D=0
M1243 395 62 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=112970 $D=0
M1244 7 63 396 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=108340 $D=0
M1245 7 63 397 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=112970 $D=0
M1246 398 64 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=108340 $D=0
M1247 399 64 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=112970 $D=0
M1248 400 396 230 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=108340 $D=0
M1249 401 397 231 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=112970 $D=0
M1250 7 400 738 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=108340 $D=0
M1251 7 401 739 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=112970 $D=0
M1252 402 738 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=108340 $D=0
M1253 403 739 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=112970 $D=0
M1254 400 63 402 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=108340 $D=0
M1255 401 63 403 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=112970 $D=0
M1256 402 398 240 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=108340 $D=0
M1257 403 399 241 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=112970 $D=0
M1258 244 404 402 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=108340 $D=0
M1259 245 405 403 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=112970 $D=0
M1260 404 65 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=108340 $D=0
M1261 405 65 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=112970 $D=0
M1262 7 66 406 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=108340 $D=0
M1263 7 66 407 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=112970 $D=0
M1264 408 67 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=108340 $D=0
M1265 409 67 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=112970 $D=0
M1266 410 406 230 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=108340 $D=0
M1267 411 407 231 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=112970 $D=0
M1268 7 410 740 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=108340 $D=0
M1269 7 411 741 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=112970 $D=0
M1270 412 740 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=108340 $D=0
M1271 413 741 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=112970 $D=0
M1272 410 66 412 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=108340 $D=0
M1273 411 66 413 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=112970 $D=0
M1274 412 408 240 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=108340 $D=0
M1275 413 409 241 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=112970 $D=0
M1276 244 414 412 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=108340 $D=0
M1277 245 415 413 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=112970 $D=0
M1278 414 68 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=108340 $D=0
M1279 415 68 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=112970 $D=0
M1280 7 69 416 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=108340 $D=0
M1281 7 69 417 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=112970 $D=0
M1282 418 70 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=108340 $D=0
M1283 419 70 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=112970 $D=0
M1284 420 416 230 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=108340 $D=0
M1285 421 417 231 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=112970 $D=0
M1286 7 420 742 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=108340 $D=0
M1287 7 421 743 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=112970 $D=0
M1288 422 742 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=108340 $D=0
M1289 423 743 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=112970 $D=0
M1290 420 69 422 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=108340 $D=0
M1291 421 69 423 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=112970 $D=0
M1292 422 418 240 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=108340 $D=0
M1293 423 419 241 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=112970 $D=0
M1294 244 424 422 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=108340 $D=0
M1295 245 425 423 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=112970 $D=0
M1296 424 71 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=108340 $D=0
M1297 425 71 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=112970 $D=0
M1298 7 72 426 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=108340 $D=0
M1299 7 72 427 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=112970 $D=0
M1300 428 73 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=108340 $D=0
M1301 429 73 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=112970 $D=0
M1302 430 426 230 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=108340 $D=0
M1303 431 427 231 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=112970 $D=0
M1304 7 430 744 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=108340 $D=0
M1305 7 431 745 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=112970 $D=0
M1306 432 744 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=108340 $D=0
M1307 433 745 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=112970 $D=0
M1308 430 72 432 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=108340 $D=0
M1309 431 72 433 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=112970 $D=0
M1310 432 428 240 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=108340 $D=0
M1311 433 429 241 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=112970 $D=0
M1312 244 434 432 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=108340 $D=0
M1313 245 435 433 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=112970 $D=0
M1314 434 74 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=108340 $D=0
M1315 435 74 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=112970 $D=0
M1316 7 75 436 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=108340 $D=0
M1317 7 75 437 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=112970 $D=0
M1318 438 76 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=108340 $D=0
M1319 439 76 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=112970 $D=0
M1320 440 436 230 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=108340 $D=0
M1321 441 437 231 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=112970 $D=0
M1322 7 440 746 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=108340 $D=0
M1323 7 441 747 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=112970 $D=0
M1324 442 746 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=108340 $D=0
M1325 443 747 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=112970 $D=0
M1326 440 75 442 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=108340 $D=0
M1327 441 75 443 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=112970 $D=0
M1328 442 438 240 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=108340 $D=0
M1329 443 439 241 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=112970 $D=0
M1330 244 444 442 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=108340 $D=0
M1331 245 445 443 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=112970 $D=0
M1332 444 77 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=108340 $D=0
M1333 445 77 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=112970 $D=0
M1334 7 78 446 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=108340 $D=0
M1335 7 78 447 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=112970 $D=0
M1336 448 79 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=108340 $D=0
M1337 449 79 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=112970 $D=0
M1338 450 446 230 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=108340 $D=0
M1339 451 447 231 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=112970 $D=0
M1340 7 450 748 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=108340 $D=0
M1341 7 451 749 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=112970 $D=0
M1342 452 748 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=108340 $D=0
M1343 453 749 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=112970 $D=0
M1344 450 78 452 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=108340 $D=0
M1345 451 78 453 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=112970 $D=0
M1346 452 448 240 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=108340 $D=0
M1347 453 449 241 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=112970 $D=0
M1348 244 454 452 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=108340 $D=0
M1349 245 455 453 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=112970 $D=0
M1350 454 80 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=108340 $D=0
M1351 455 80 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=112970 $D=0
M1352 7 81 456 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=108340 $D=0
M1353 7 81 457 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=112970 $D=0
M1354 458 82 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=108340 $D=0
M1355 459 82 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=112970 $D=0
M1356 460 456 230 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=108340 $D=0
M1357 461 457 231 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=112970 $D=0
M1358 7 460 750 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=108340 $D=0
M1359 7 461 751 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=112970 $D=0
M1360 462 750 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=108340 $D=0
M1361 463 751 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=112970 $D=0
M1362 460 81 462 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=108340 $D=0
M1363 461 81 463 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=112970 $D=0
M1364 462 458 240 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=108340 $D=0
M1365 463 459 241 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=112970 $D=0
M1366 244 464 462 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=108340 $D=0
M1367 245 465 463 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=112970 $D=0
M1368 464 83 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=108340 $D=0
M1369 465 83 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=112970 $D=0
M1370 7 84 466 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=108340 $D=0
M1371 7 84 467 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=112970 $D=0
M1372 468 85 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=108340 $D=0
M1373 469 85 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=112970 $D=0
M1374 470 466 230 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=108340 $D=0
M1375 471 467 231 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=112970 $D=0
M1376 7 470 752 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=108340 $D=0
M1377 7 471 753 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=112970 $D=0
M1378 472 752 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=108340 $D=0
M1379 473 753 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=112970 $D=0
M1380 470 84 472 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=108340 $D=0
M1381 471 84 473 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=112970 $D=0
M1382 472 468 240 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=108340 $D=0
M1383 473 469 241 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=112970 $D=0
M1384 244 474 472 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=108340 $D=0
M1385 245 475 473 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=112970 $D=0
M1386 474 86 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=108340 $D=0
M1387 475 86 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=112970 $D=0
M1388 7 87 476 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=108340 $D=0
M1389 7 87 477 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=112970 $D=0
M1390 478 88 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=108340 $D=0
M1391 479 88 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=112970 $D=0
M1392 480 476 230 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=108340 $D=0
M1393 481 477 231 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=112970 $D=0
M1394 7 480 754 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=108340 $D=0
M1395 7 481 755 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=112970 $D=0
M1396 482 754 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=108340 $D=0
M1397 483 755 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=112970 $D=0
M1398 480 87 482 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=108340 $D=0
M1399 481 87 483 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=112970 $D=0
M1400 482 478 240 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=108340 $D=0
M1401 483 479 241 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=112970 $D=0
M1402 244 484 482 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=108340 $D=0
M1403 245 485 483 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=112970 $D=0
M1404 484 89 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=108340 $D=0
M1405 485 89 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=112970 $D=0
M1406 7 90 486 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=108340 $D=0
M1407 7 90 487 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=112970 $D=0
M1408 488 91 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=108340 $D=0
M1409 489 91 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=112970 $D=0
M1410 490 486 230 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=108340 $D=0
M1411 491 487 231 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=112970 $D=0
M1412 7 490 756 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=108340 $D=0
M1413 7 491 757 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=112970 $D=0
M1414 492 756 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=108340 $D=0
M1415 493 757 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=112970 $D=0
M1416 490 90 492 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=108340 $D=0
M1417 491 90 493 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=112970 $D=0
M1418 492 488 240 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=108340 $D=0
M1419 493 489 241 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=112970 $D=0
M1420 244 494 492 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=108340 $D=0
M1421 245 495 493 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=112970 $D=0
M1422 494 92 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=108340 $D=0
M1423 495 92 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=112970 $D=0
M1424 7 93 496 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=108340 $D=0
M1425 7 93 497 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=112970 $D=0
M1426 498 94 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=108340 $D=0
M1427 499 94 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=112970 $D=0
M1428 500 496 230 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=108340 $D=0
M1429 501 497 231 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=112970 $D=0
M1430 7 500 758 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=108340 $D=0
M1431 7 501 759 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=112970 $D=0
M1432 502 758 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=108340 $D=0
M1433 503 759 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=112970 $D=0
M1434 500 93 502 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=108340 $D=0
M1435 501 93 503 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=112970 $D=0
M1436 502 498 240 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=108340 $D=0
M1437 503 499 241 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=112970 $D=0
M1438 244 504 502 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=108340 $D=0
M1439 245 505 503 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=112970 $D=0
M1440 504 95 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=108340 $D=0
M1441 505 95 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=112970 $D=0
M1442 7 96 506 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=108340 $D=0
M1443 7 96 507 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=112970 $D=0
M1444 508 97 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=108340 $D=0
M1445 509 97 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=112970 $D=0
M1446 510 506 230 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=108340 $D=0
M1447 511 507 231 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=112970 $D=0
M1448 7 510 760 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=108340 $D=0
M1449 7 511 761 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=112970 $D=0
M1450 512 760 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=108340 $D=0
M1451 513 761 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=112970 $D=0
M1452 510 96 512 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=108340 $D=0
M1453 511 96 513 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=112970 $D=0
M1454 512 508 240 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=108340 $D=0
M1455 513 509 241 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=112970 $D=0
M1456 244 514 512 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=108340 $D=0
M1457 245 515 513 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=112970 $D=0
M1458 514 98 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=108340 $D=0
M1459 515 98 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=112970 $D=0
M1460 7 99 516 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=108340 $D=0
M1461 7 99 517 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=112970 $D=0
M1462 518 100 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=108340 $D=0
M1463 519 100 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=112970 $D=0
M1464 520 516 230 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=108340 $D=0
M1465 521 517 231 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=112970 $D=0
M1466 7 520 762 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=108340 $D=0
M1467 7 521 763 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=112970 $D=0
M1468 522 762 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=108340 $D=0
M1469 523 763 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=112970 $D=0
M1470 520 99 522 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=108340 $D=0
M1471 521 99 523 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=112970 $D=0
M1472 522 518 240 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=108340 $D=0
M1473 523 519 241 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=112970 $D=0
M1474 244 524 522 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=108340 $D=0
M1475 245 525 523 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=112970 $D=0
M1476 524 101 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=108340 $D=0
M1477 525 101 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=112970 $D=0
M1478 7 102 526 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=108340 $D=0
M1479 7 102 527 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=112970 $D=0
M1480 528 103 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=108340 $D=0
M1481 529 103 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=112970 $D=0
M1482 530 526 230 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=108340 $D=0
M1483 531 527 231 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=112970 $D=0
M1484 7 530 764 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=108340 $D=0
M1485 7 531 765 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=112970 $D=0
M1486 532 764 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=108340 $D=0
M1487 533 765 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=112970 $D=0
M1488 530 102 532 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=108340 $D=0
M1489 531 102 533 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=112970 $D=0
M1490 532 528 240 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=108340 $D=0
M1491 533 529 241 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=112970 $D=0
M1492 244 534 532 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=108340 $D=0
M1493 245 535 533 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=112970 $D=0
M1494 534 104 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=108340 $D=0
M1495 535 104 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=112970 $D=0
M1496 7 105 536 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=108340 $D=0
M1497 7 105 537 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=112970 $D=0
M1498 538 106 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=108340 $D=0
M1499 539 106 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=112970 $D=0
M1500 540 536 230 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=108340 $D=0
M1501 541 537 231 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=112970 $D=0
M1502 7 540 766 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=108340 $D=0
M1503 7 541 767 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=112970 $D=0
M1504 542 766 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=108340 $D=0
M1505 543 767 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=112970 $D=0
M1506 540 105 542 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=108340 $D=0
M1507 541 105 543 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=112970 $D=0
M1508 542 538 240 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=108340 $D=0
M1509 543 539 241 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=112970 $D=0
M1510 244 544 542 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=108340 $D=0
M1511 245 545 543 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=112970 $D=0
M1512 544 107 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=108340 $D=0
M1513 545 107 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=112970 $D=0
M1514 7 108 546 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=108340 $D=0
M1515 7 108 547 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=112970 $D=0
M1516 548 109 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=108340 $D=0
M1517 549 109 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=112970 $D=0
M1518 4 548 240 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=108340 $D=0
M1519 4 549 241 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=112970 $D=0
M1520 244 546 4 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=108340 $D=0
M1521 245 547 4 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=112970 $D=0
M1522 7 552 550 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=108340 $D=0
M1523 7 553 551 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=112970 $D=0
M1524 552 110 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=108340 $D=0
M1525 553 110 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=112970 $D=0
M1526 768 240 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=108340 $D=0
M1527 769 241 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=112970 $D=0
M1528 554 552 768 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=108340 $D=0
M1529 555 553 769 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=112970 $D=0
M1530 7 554 556 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=108340 $D=0
M1531 7 555 557 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=112970 $D=0
M1532 770 556 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=108340 $D=0
M1533 771 557 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=112970 $D=0
M1534 554 550 770 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=108340 $D=0
M1535 555 551 771 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=112970 $D=0
M1536 7 560 558 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=108340 $D=0
M1537 7 561 559 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=112970 $D=0
M1538 560 110 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=108340 $D=0
M1539 561 110 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=112970 $D=0
M1540 772 244 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=108340 $D=0
M1541 773 245 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=112970 $D=0
M1542 562 560 772 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=108340 $D=0
M1543 563 561 773 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=112970 $D=0
M1544 7 562 111 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=108340 $D=0
M1545 7 563 112 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=112970 $D=0
M1546 774 111 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=108340 $D=0
M1547 775 112 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=112970 $D=0
M1548 562 558 774 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=108340 $D=0
M1549 563 559 775 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=112970 $D=0
M1550 564 113 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=108340 $D=0
M1551 565 113 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=112970 $D=0
M1552 566 113 556 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=108340 $D=0
M1553 567 113 557 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=112970 $D=0
M1554 114 564 566 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=108340 $D=0
M1555 115 565 567 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=112970 $D=0
M1556 568 116 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=108340 $D=0
M1557 569 116 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=112970 $D=0
M1558 570 116 111 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=108340 $D=0
M1559 571 116 112 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=112970 $D=0
M1560 776 568 570 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=108340 $D=0
M1561 777 569 571 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=112970 $D=0
M1562 7 111 776 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=108340 $D=0
M1563 7 112 777 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=112970 $D=0
M1564 572 118 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=108340 $D=0
M1565 573 118 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=112970 $D=0
M1566 574 118 570 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=108340 $D=0
M1567 575 118 571 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=112970 $D=0
M1568 9 572 574 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=108340 $D=0
M1569 10 573 575 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=112970 $D=0
M1570 577 576 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=108340 $D=0
M1571 578 120 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=112970 $D=0
M1572 7 581 579 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=108340 $D=0
M1573 7 582 580 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=112970 $D=0
M1574 583 566 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=108340 $D=0
M1575 584 567 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=112970 $D=0
M1576 581 566 576 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=108340 $D=0
M1577 582 567 120 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=112970 $D=0
M1578 577 583 581 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=108340 $D=0
M1579 578 584 582 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=112970 $D=0
M1580 585 579 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=108340 $D=0
M1581 586 580 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=112970 $D=0
M1582 124 579 574 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=108340 $D=0
M1583 576 580 575 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=112970 $D=0
M1584 566 585 124 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=108340 $D=0
M1585 567 586 576 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=112970 $D=0
M1586 587 124 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=108340 $D=0
M1587 588 576 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=112970 $D=0
M1588 589 579 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=108340 $D=0
M1589 590 580 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=112970 $D=0
M1590 591 579 587 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=108340 $D=0
M1591 592 580 588 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=112970 $D=0
M1592 574 589 591 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=108340 $D=0
M1593 575 590 592 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=112970 $D=0
M1594 788 566 7 7 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=107980 $D=0
M1595 789 567 7 7 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=112610 $D=0
M1596 593 574 788 7 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=107980 $D=0
M1597 594 575 789 7 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=112610 $D=0
M1598 595 591 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=108340 $D=0
M1599 596 592 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=112970 $D=0
M1600 597 566 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=108340 $D=0
M1601 598 567 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=112970 $D=0
M1602 7 574 597 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=108340 $D=0
M1603 7 575 598 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=112970 $D=0
M1604 599 566 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=108340 $D=0
M1605 600 567 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=112970 $D=0
M1606 7 574 599 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=108340 $D=0
M1607 7 575 600 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=112970 $D=0
M1608 790 566 7 7 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=108160 $D=0
M1609 791 567 7 7 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=112790 $D=0
M1610 603 574 790 7 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=108160 $D=0
M1611 604 575 791 7 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=112790 $D=0
M1612 7 599 603 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=108340 $D=0
M1613 7 600 604 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=112970 $D=0
M1614 605 126 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=108340 $D=0
M1615 606 126 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=112970 $D=0
M1616 607 126 593 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=108340 $D=0
M1617 608 126 594 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=112970 $D=0
M1618 597 605 607 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=108340 $D=0
M1619 598 606 608 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=112970 $D=0
M1620 609 126 595 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=108340 $D=0
M1621 610 126 596 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=112970 $D=0
M1622 603 605 609 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=108340 $D=0
M1623 604 606 610 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=112970 $D=0
M1624 611 127 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=108340 $D=0
M1625 612 127 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=112970 $D=0
M1626 613 127 609 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=108340 $D=0
M1627 614 127 610 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=112970 $D=0
M1628 607 611 613 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=108340 $D=0
M1629 608 612 614 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=112970 $D=0
M1630 11 613 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=108340 $D=0
M1631 12 614 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=112970 $D=0
M1632 615 128 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=108340 $D=0
M1633 616 128 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=112970 $D=0
M1634 617 128 129 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=108340 $D=0
M1635 618 128 130 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=112970 $D=0
M1636 131 615 617 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=108340 $D=0
M1637 132 616 618 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=112970 $D=0
M1638 619 128 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=108340 $D=0
M1639 620 128 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=112970 $D=0
M1640 621 128 133 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=108340 $D=0
M1641 622 128 134 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=112970 $D=0
M1642 135 619 621 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=108340 $D=0
M1643 136 620 622 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=112970 $D=0
M1644 623 128 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=108340 $D=0
M1645 624 128 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=112970 $D=0
M1646 625 128 137 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=108340 $D=0
M1647 626 128 138 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=112970 $D=0
M1648 117 623 625 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=108340 $D=0
M1649 123 624 626 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=112970 $D=0
M1650 627 128 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=108340 $D=0
M1651 628 128 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=112970 $D=0
M1652 629 128 139 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=108340 $D=0
M1653 630 128 4 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=112970 $D=0
M1654 119 627 629 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=108340 $D=0
M1655 140 628 630 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=112970 $D=0
M1656 631 128 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=108340 $D=0
M1657 632 128 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=112970 $D=0
M1658 633 128 4 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=108340 $D=0
M1659 634 128 4 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=112970 $D=0
M1660 141 631 633 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=108340 $D=0
M1661 142 632 634 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=112970 $D=0
M1662 7 566 778 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=108340 $D=0
M1663 7 567 779 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=112970 $D=0
M1664 132 778 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=108340 $D=0
M1665 129 779 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=112970 $D=0
M1666 635 143 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=108340 $D=0
M1667 636 143 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=112970 $D=0
M1668 144 143 132 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=108340 $D=0
M1669 145 143 129 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=112970 $D=0
M1670 617 635 144 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=108340 $D=0
M1671 618 636 145 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=112970 $D=0
M1672 637 146 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=108340 $D=0
M1673 638 146 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=112970 $D=0
M1674 125 146 144 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=108340 $D=0
M1675 147 146 145 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=112970 $D=0
M1676 621 637 125 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=108340 $D=0
M1677 622 638 147 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=112970 $D=0
M1678 639 148 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=108340 $D=0
M1679 640 148 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=112970 $D=0
M1680 121 148 125 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=108340 $D=0
M1681 122 148 147 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=112970 $D=0
M1682 625 639 121 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=108340 $D=0
M1683 626 640 122 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=112970 $D=0
M1684 641 149 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=108340 $D=0
M1685 642 149 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=112970 $D=0
M1686 150 149 121 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=108340 $D=0
M1687 151 149 122 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=112970 $D=0
M1688 629 641 150 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=108340 $D=0
M1689 630 642 151 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=112970 $D=0
M1690 643 152 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=108340 $D=0
M1691 644 152 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=112970 $D=0
M1692 216 152 150 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=108340 $D=0
M1693 217 152 151 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=112970 $D=0
M1694 633 643 216 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=108340 $D=0
M1695 634 644 217 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=112970 $D=0
M1696 645 153 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=108340 $D=0
M1697 646 153 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=112970 $D=0
M1698 647 153 111 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=108340 $D=0
M1699 648 153 112 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=112970 $D=0
M1700 9 645 647 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=108340 $D=0
M1701 10 646 648 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=112970 $D=0
M1702 649 556 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=108340 $D=0
M1703 650 557 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=112970 $D=0
M1704 7 647 649 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=108340 $D=0
M1705 7 648 650 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=112970 $D=0
M1706 792 556 7 7 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=108160 $D=0
M1707 793 557 7 7 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=112790 $D=0
M1708 653 647 792 7 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=108160 $D=0
M1709 654 648 793 7 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=112790 $D=0
M1710 7 649 653 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=108340 $D=0
M1711 7 650 654 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=112970 $D=0
M1712 780 154 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=108340 $D=0
M1713 781 655 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=112970 $D=0
M1714 7 653 780 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=108340 $D=0
M1715 7 654 781 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=112970 $D=0
M1716 655 780 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=108340 $D=0
M1717 155 781 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=112970 $D=0
M1718 794 556 7 7 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=107980 $D=0
M1719 795 557 7 7 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=112610 $D=0
M1720 656 658 794 7 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=107980 $D=0
M1721 657 659 795 7 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=112610 $D=0
M1722 658 647 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=108340 $D=0
M1723 659 648 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=112970 $D=0
M1724 660 656 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=108340 $D=0
M1725 661 657 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=112970 $D=0
M1726 7 154 660 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=108340 $D=0
M1727 7 655 661 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=112970 $D=0
M1728 663 156 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=108340 $D=0
M1729 664 662 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=112970 $D=0
M1730 662 660 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=108340 $D=0
M1731 157 661 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=112970 $D=0
M1732 7 663 662 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=108340 $D=0
M1733 7 664 157 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=112970 $D=0
M1734 666 665 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=108340 $D=0
M1735 667 158 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=112970 $D=0
M1736 7 670 668 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=108340 $D=0
M1737 7 671 669 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=112970 $D=0
M1738 672 114 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=108340 $D=0
M1739 673 115 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=112970 $D=0
M1740 670 114 665 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=108340 $D=0
M1741 671 115 158 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=112970 $D=0
M1742 666 672 670 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=108340 $D=0
M1743 667 673 671 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=112970 $D=0
M1744 674 668 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=108340 $D=0
M1745 675 669 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=112970 $D=0
M1746 159 668 4 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=108340 $D=0
M1747 665 669 4 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=112970 $D=0
M1748 114 674 159 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=108340 $D=0
M1749 115 675 665 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=112970 $D=0
M1750 676 159 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=108340 $D=0
M1751 677 665 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=112970 $D=0
M1752 678 668 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=108340 $D=0
M1753 679 669 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=112970 $D=0
M1754 218 668 676 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=108340 $D=0
M1755 219 669 677 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=112970 $D=0
M1756 4 678 218 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=108340 $D=0
M1757 4 679 219 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=112970 $D=0
M1758 680 160 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=108340 $D=0
M1759 681 160 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=112970 $D=0
M1760 682 160 218 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=108340 $D=0
M1761 683 160 219 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=112970 $D=0
M1762 11 680 682 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=108340 $D=0
M1763 12 681 683 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=112970 $D=0
M1764 684 161 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=108340 $D=0
M1765 685 161 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=112970 $D=0
M1766 686 161 682 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=108340 $D=0
M1767 687 161 683 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=112970 $D=0
M1768 4 684 686 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=108340 $D=0
M1769 4 685 687 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=112970 $D=0
M1770 688 110 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=108340 $D=0
M1771 689 110 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=112970 $D=0
M1772 7 688 690 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=108340 $D=0
M1773 7 689 691 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=112970 $D=0
M1774 692 110 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=108340 $D=0
M1775 693 110 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=112970 $D=0
M1776 694 690 686 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=108340 $D=0
M1777 695 691 687 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=112970 $D=0
M1778 7 694 782 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=108340 $D=0
M1779 7 695 783 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=112970 $D=0
M1780 696 782 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=108340 $D=0
M1781 697 783 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=112970 $D=0
M1782 694 688 696 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=108340 $D=0
M1783 695 689 697 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=112970 $D=0
M1784 698 692 696 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=108340 $D=0
M1785 699 693 697 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=112970 $D=0
M1786 7 702 700 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=108340 $D=0
M1787 7 703 701 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=112970 $D=0
M1788 702 110 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=108340 $D=0
M1789 703 110 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=112970 $D=0
M1790 784 698 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=108340 $D=0
M1791 785 699 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=112970 $D=0
M1792 704 702 784 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=108340 $D=0
M1793 705 703 785 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=112970 $D=0
M1794 7 704 114 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=108340 $D=0
M1795 7 705 115 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=112970 $D=0
M1796 786 114 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=108340 $D=0
M1797 787 115 7 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=112970 $D=0
M1798 704 700 786 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=108340 $D=0
M1799 705 701 787 7 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=112970 $D=0
.ENDS
***************************************
.SUBCKT ICV_28 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163
** N=813 EP=163 IP=1514 FDC=1800
M0 198 1 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=97830 $D=1
M1 199 1 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=102460 $D=1
M2 200 198 2 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=97830 $D=1
M3 201 199 3 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=102460 $D=1
M4 5 1 200 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=97830 $D=1
M5 5 1 201 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=102460 $D=1
M6 202 198 4 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=97830 $D=1
M7 203 199 4 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=102460 $D=1
M8 2 1 202 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=97830 $D=1
M9 3 1 203 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=102460 $D=1
M10 204 198 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=97830 $D=1
M11 205 199 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=102460 $D=1
M12 2 1 204 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=97830 $D=1
M13 3 1 205 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=102460 $D=1
M14 208 206 204 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=97830 $D=1
M15 209 207 205 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=102460 $D=1
M16 206 6 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=97830 $D=1
M17 207 6 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=102460 $D=1
M18 210 206 202 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=97830 $D=1
M19 211 207 203 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=102460 $D=1
M20 200 6 210 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=97830 $D=1
M21 201 6 211 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=102460 $D=1
M22 212 7 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=97830 $D=1
M23 213 7 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=102460 $D=1
M24 214 212 210 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=97830 $D=1
M25 215 213 211 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=102460 $D=1
M26 208 7 214 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=97830 $D=1
M27 209 7 215 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=102460 $D=1
M28 216 9 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=97830 $D=1
M29 217 9 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=102460 $D=1
M30 218 216 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=97830 $D=1
M31 219 217 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=102460 $D=1
M32 10 9 218 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=97830 $D=1
M33 11 9 219 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=102460 $D=1
M34 220 216 12 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=97830 $D=1
M35 221 217 13 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=102460 $D=1
M36 222 9 220 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=97830 $D=1
M37 223 9 221 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=102460 $D=1
M38 226 216 224 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=97830 $D=1
M39 227 217 225 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=102460 $D=1
M40 214 9 226 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=97830 $D=1
M41 215 9 227 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=102460 $D=1
M42 230 228 226 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=97830 $D=1
M43 231 229 227 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=102460 $D=1
M44 228 14 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=97830 $D=1
M45 229 14 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=102460 $D=1
M46 232 228 220 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=97830 $D=1
M47 233 229 221 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=102460 $D=1
M48 218 14 232 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=97830 $D=1
M49 219 14 233 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=102460 $D=1
M50 234 15 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=97830 $D=1
M51 235 15 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=102460 $D=1
M52 236 234 232 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=97830 $D=1
M53 237 235 233 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=102460 $D=1
M54 230 15 236 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=97830 $D=1
M55 231 15 237 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=102460 $D=1
M56 5 16 238 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=97830 $D=1
M57 5 16 239 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=102460 $D=1
M58 240 17 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=97830 $D=1
M59 241 17 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=102460 $D=1
M60 242 16 236 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=97830 $D=1
M61 243 16 237 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=102460 $D=1
M62 5 242 712 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=97830 $D=1
M63 5 243 713 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=102460 $D=1
M64 244 712 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=97830 $D=1
M65 245 713 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=102460 $D=1
M66 242 238 244 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=97830 $D=1
M67 243 239 245 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=102460 $D=1
M68 244 17 246 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=97830 $D=1
M69 245 17 247 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=102460 $D=1
M70 250 18 244 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=97830 $D=1
M71 251 18 245 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=102460 $D=1
M72 248 18 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=97830 $D=1
M73 249 18 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=102460 $D=1
M74 5 19 252 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=97830 $D=1
M75 5 19 253 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=102460 $D=1
M76 254 20 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=97830 $D=1
M77 255 20 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=102460 $D=1
M78 256 19 236 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=97830 $D=1
M79 257 19 237 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=102460 $D=1
M80 5 256 714 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=97830 $D=1
M81 5 257 715 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=102460 $D=1
M82 258 714 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=97830 $D=1
M83 259 715 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=102460 $D=1
M84 256 252 258 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=97830 $D=1
M85 257 253 259 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=102460 $D=1
M86 258 20 246 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=97830 $D=1
M87 259 20 247 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=102460 $D=1
M88 250 21 258 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=97830 $D=1
M89 251 21 259 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=102460 $D=1
M90 260 21 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=97830 $D=1
M91 261 21 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=102460 $D=1
M92 5 22 262 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=97830 $D=1
M93 5 22 263 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=102460 $D=1
M94 264 23 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=97830 $D=1
M95 265 23 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=102460 $D=1
M96 266 22 236 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=97830 $D=1
M97 267 22 237 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=102460 $D=1
M98 5 266 716 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=97830 $D=1
M99 5 267 717 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=102460 $D=1
M100 268 716 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=97830 $D=1
M101 269 717 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=102460 $D=1
M102 266 262 268 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=97830 $D=1
M103 267 263 269 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=102460 $D=1
M104 268 23 246 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=97830 $D=1
M105 269 23 247 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=102460 $D=1
M106 250 24 268 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=97830 $D=1
M107 251 24 269 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=102460 $D=1
M108 270 24 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=97830 $D=1
M109 271 24 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=102460 $D=1
M110 5 25 272 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=97830 $D=1
M111 5 25 273 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=102460 $D=1
M112 274 26 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=97830 $D=1
M113 275 26 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=102460 $D=1
M114 276 25 236 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=97830 $D=1
M115 277 25 237 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=102460 $D=1
M116 5 276 718 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=97830 $D=1
M117 5 277 719 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=102460 $D=1
M118 278 718 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=97830 $D=1
M119 279 719 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=102460 $D=1
M120 276 272 278 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=97830 $D=1
M121 277 273 279 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=102460 $D=1
M122 278 26 246 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=97830 $D=1
M123 279 26 247 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=102460 $D=1
M124 250 27 278 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=97830 $D=1
M125 251 27 279 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=102460 $D=1
M126 280 27 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=97830 $D=1
M127 281 27 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=102460 $D=1
M128 5 28 282 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=97830 $D=1
M129 5 28 283 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=102460 $D=1
M130 284 29 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=97830 $D=1
M131 285 29 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=102460 $D=1
M132 286 28 236 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=97830 $D=1
M133 287 28 237 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=102460 $D=1
M134 5 286 720 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=97830 $D=1
M135 5 287 721 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=102460 $D=1
M136 288 720 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=97830 $D=1
M137 289 721 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=102460 $D=1
M138 286 282 288 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=97830 $D=1
M139 287 283 289 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=102460 $D=1
M140 288 29 246 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=97830 $D=1
M141 289 29 247 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=102460 $D=1
M142 250 30 288 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=97830 $D=1
M143 251 30 289 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=102460 $D=1
M144 290 30 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=97830 $D=1
M145 291 30 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=102460 $D=1
M146 5 31 292 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=97830 $D=1
M147 5 31 293 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=102460 $D=1
M148 294 32 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=97830 $D=1
M149 295 32 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=102460 $D=1
M150 296 31 236 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=97830 $D=1
M151 297 31 237 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=102460 $D=1
M152 5 296 722 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=97830 $D=1
M153 5 297 723 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=102460 $D=1
M154 298 722 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=97830 $D=1
M155 299 723 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=102460 $D=1
M156 296 292 298 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=97830 $D=1
M157 297 293 299 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=102460 $D=1
M158 298 32 246 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=97830 $D=1
M159 299 32 247 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=102460 $D=1
M160 250 33 298 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=97830 $D=1
M161 251 33 299 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=102460 $D=1
M162 300 33 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=97830 $D=1
M163 301 33 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=102460 $D=1
M164 5 34 302 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=97830 $D=1
M165 5 34 303 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=102460 $D=1
M166 304 35 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=97830 $D=1
M167 305 35 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=102460 $D=1
M168 306 34 236 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=97830 $D=1
M169 307 34 237 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=102460 $D=1
M170 5 306 724 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=97830 $D=1
M171 5 307 725 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=102460 $D=1
M172 308 724 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=97830 $D=1
M173 309 725 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=102460 $D=1
M174 306 302 308 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=97830 $D=1
M175 307 303 309 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=102460 $D=1
M176 308 35 246 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=97830 $D=1
M177 309 35 247 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=102460 $D=1
M178 250 36 308 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=97830 $D=1
M179 251 36 309 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=102460 $D=1
M180 310 36 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=97830 $D=1
M181 311 36 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=102460 $D=1
M182 5 37 312 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=97830 $D=1
M183 5 37 313 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=102460 $D=1
M184 314 38 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=97830 $D=1
M185 315 38 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=102460 $D=1
M186 316 37 236 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=97830 $D=1
M187 317 37 237 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=102460 $D=1
M188 5 316 726 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=97830 $D=1
M189 5 317 727 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=102460 $D=1
M190 318 726 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=97830 $D=1
M191 319 727 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=102460 $D=1
M192 316 312 318 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=97830 $D=1
M193 317 313 319 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=102460 $D=1
M194 318 38 246 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=97830 $D=1
M195 319 38 247 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=102460 $D=1
M196 250 39 318 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=97830 $D=1
M197 251 39 319 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=102460 $D=1
M198 320 39 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=97830 $D=1
M199 321 39 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=102460 $D=1
M200 5 40 322 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=97830 $D=1
M201 5 40 323 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=102460 $D=1
M202 324 41 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=97830 $D=1
M203 325 41 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=102460 $D=1
M204 326 40 236 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=97830 $D=1
M205 327 40 237 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=102460 $D=1
M206 5 326 728 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=97830 $D=1
M207 5 327 729 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=102460 $D=1
M208 328 728 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=97830 $D=1
M209 329 729 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=102460 $D=1
M210 326 322 328 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=97830 $D=1
M211 327 323 329 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=102460 $D=1
M212 328 41 246 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=97830 $D=1
M213 329 41 247 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=102460 $D=1
M214 250 42 328 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=97830 $D=1
M215 251 42 329 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=102460 $D=1
M216 330 42 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=97830 $D=1
M217 331 42 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=102460 $D=1
M218 5 43 332 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=97830 $D=1
M219 5 43 333 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=102460 $D=1
M220 334 44 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=97830 $D=1
M221 335 44 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=102460 $D=1
M222 336 43 236 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=97830 $D=1
M223 337 43 237 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=102460 $D=1
M224 5 336 730 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=97830 $D=1
M225 5 337 731 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=102460 $D=1
M226 338 730 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=97830 $D=1
M227 339 731 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=102460 $D=1
M228 336 332 338 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=97830 $D=1
M229 337 333 339 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=102460 $D=1
M230 338 44 246 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=97830 $D=1
M231 339 44 247 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=102460 $D=1
M232 250 45 338 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=97830 $D=1
M233 251 45 339 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=102460 $D=1
M234 340 45 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=97830 $D=1
M235 341 45 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=102460 $D=1
M236 5 46 342 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=97830 $D=1
M237 5 46 343 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=102460 $D=1
M238 344 47 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=97830 $D=1
M239 345 47 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=102460 $D=1
M240 346 46 236 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=97830 $D=1
M241 347 46 237 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=102460 $D=1
M242 5 346 732 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=97830 $D=1
M243 5 347 733 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=102460 $D=1
M244 348 732 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=97830 $D=1
M245 349 733 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=102460 $D=1
M246 346 342 348 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=97830 $D=1
M247 347 343 349 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=102460 $D=1
M248 348 47 246 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=97830 $D=1
M249 349 47 247 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=102460 $D=1
M250 250 48 348 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=97830 $D=1
M251 251 48 349 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=102460 $D=1
M252 350 48 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=97830 $D=1
M253 351 48 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=102460 $D=1
M254 5 49 352 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=97830 $D=1
M255 5 49 353 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=102460 $D=1
M256 354 50 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=97830 $D=1
M257 355 50 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=102460 $D=1
M258 356 49 236 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=97830 $D=1
M259 357 49 237 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=102460 $D=1
M260 5 356 734 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=97830 $D=1
M261 5 357 735 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=102460 $D=1
M262 358 734 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=97830 $D=1
M263 359 735 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=102460 $D=1
M264 356 352 358 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=97830 $D=1
M265 357 353 359 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=102460 $D=1
M266 358 50 246 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=97830 $D=1
M267 359 50 247 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=102460 $D=1
M268 250 51 358 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=97830 $D=1
M269 251 51 359 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=102460 $D=1
M270 360 51 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=97830 $D=1
M271 361 51 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=102460 $D=1
M272 5 52 362 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=97830 $D=1
M273 5 52 363 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=102460 $D=1
M274 364 53 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=97830 $D=1
M275 365 53 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=102460 $D=1
M276 366 52 236 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=97830 $D=1
M277 367 52 237 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=102460 $D=1
M278 5 366 736 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=97830 $D=1
M279 5 367 737 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=102460 $D=1
M280 368 736 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=97830 $D=1
M281 369 737 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=102460 $D=1
M282 366 362 368 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=97830 $D=1
M283 367 363 369 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=102460 $D=1
M284 368 53 246 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=97830 $D=1
M285 369 53 247 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=102460 $D=1
M286 250 54 368 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=97830 $D=1
M287 251 54 369 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=102460 $D=1
M288 370 54 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=97830 $D=1
M289 371 54 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=102460 $D=1
M290 5 55 372 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=97830 $D=1
M291 5 55 373 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=102460 $D=1
M292 374 56 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=97830 $D=1
M293 375 56 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=102460 $D=1
M294 376 55 236 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=97830 $D=1
M295 377 55 237 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=102460 $D=1
M296 5 376 738 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=97830 $D=1
M297 5 377 739 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=102460 $D=1
M298 378 738 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=97830 $D=1
M299 379 739 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=102460 $D=1
M300 376 372 378 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=97830 $D=1
M301 377 373 379 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=102460 $D=1
M302 378 56 246 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=97830 $D=1
M303 379 56 247 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=102460 $D=1
M304 250 57 378 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=97830 $D=1
M305 251 57 379 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=102460 $D=1
M306 380 57 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=97830 $D=1
M307 381 57 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=102460 $D=1
M308 5 58 382 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=97830 $D=1
M309 5 58 383 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=102460 $D=1
M310 384 59 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=97830 $D=1
M311 385 59 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=102460 $D=1
M312 386 58 236 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=97830 $D=1
M313 387 58 237 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=102460 $D=1
M314 5 386 740 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=97830 $D=1
M315 5 387 741 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=102460 $D=1
M316 388 740 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=97830 $D=1
M317 389 741 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=102460 $D=1
M318 386 382 388 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=97830 $D=1
M319 387 383 389 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=102460 $D=1
M320 388 59 246 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=97830 $D=1
M321 389 59 247 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=102460 $D=1
M322 250 60 388 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=97830 $D=1
M323 251 60 389 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=102460 $D=1
M324 390 60 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=97830 $D=1
M325 391 60 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=102460 $D=1
M326 5 61 392 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=97830 $D=1
M327 5 61 393 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=102460 $D=1
M328 394 62 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=97830 $D=1
M329 395 62 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=102460 $D=1
M330 396 61 236 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=97830 $D=1
M331 397 61 237 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=102460 $D=1
M332 5 396 742 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=97830 $D=1
M333 5 397 743 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=102460 $D=1
M334 398 742 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=97830 $D=1
M335 399 743 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=102460 $D=1
M336 396 392 398 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=97830 $D=1
M337 397 393 399 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=102460 $D=1
M338 398 62 246 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=97830 $D=1
M339 399 62 247 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=102460 $D=1
M340 250 63 398 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=97830 $D=1
M341 251 63 399 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=102460 $D=1
M342 400 63 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=97830 $D=1
M343 401 63 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=102460 $D=1
M344 5 64 402 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=97830 $D=1
M345 5 64 403 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=102460 $D=1
M346 404 65 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=97830 $D=1
M347 405 65 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=102460 $D=1
M348 406 64 236 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=97830 $D=1
M349 407 64 237 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=102460 $D=1
M350 5 406 744 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=97830 $D=1
M351 5 407 745 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=102460 $D=1
M352 408 744 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=97830 $D=1
M353 409 745 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=102460 $D=1
M354 406 402 408 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=97830 $D=1
M355 407 403 409 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=102460 $D=1
M356 408 65 246 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=97830 $D=1
M357 409 65 247 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=102460 $D=1
M358 250 66 408 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=97830 $D=1
M359 251 66 409 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=102460 $D=1
M360 410 66 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=97830 $D=1
M361 411 66 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=102460 $D=1
M362 5 67 412 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=97830 $D=1
M363 5 67 413 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=102460 $D=1
M364 414 68 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=97830 $D=1
M365 415 68 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=102460 $D=1
M366 416 67 236 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=97830 $D=1
M367 417 67 237 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=102460 $D=1
M368 5 416 746 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=97830 $D=1
M369 5 417 747 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=102460 $D=1
M370 418 746 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=97830 $D=1
M371 419 747 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=102460 $D=1
M372 416 412 418 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=97830 $D=1
M373 417 413 419 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=102460 $D=1
M374 418 68 246 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=97830 $D=1
M375 419 68 247 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=102460 $D=1
M376 250 69 418 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=97830 $D=1
M377 251 69 419 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=102460 $D=1
M378 420 69 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=97830 $D=1
M379 421 69 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=102460 $D=1
M380 5 70 422 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=97830 $D=1
M381 5 70 423 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=102460 $D=1
M382 424 71 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=97830 $D=1
M383 425 71 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=102460 $D=1
M384 426 70 236 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=97830 $D=1
M385 427 70 237 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=102460 $D=1
M386 5 426 748 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=97830 $D=1
M387 5 427 749 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=102460 $D=1
M388 428 748 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=97830 $D=1
M389 429 749 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=102460 $D=1
M390 426 422 428 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=97830 $D=1
M391 427 423 429 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=102460 $D=1
M392 428 71 246 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=97830 $D=1
M393 429 71 247 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=102460 $D=1
M394 250 72 428 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=97830 $D=1
M395 251 72 429 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=102460 $D=1
M396 430 72 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=97830 $D=1
M397 431 72 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=102460 $D=1
M398 5 73 432 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=97830 $D=1
M399 5 73 433 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=102460 $D=1
M400 434 74 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=97830 $D=1
M401 435 74 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=102460 $D=1
M402 436 73 236 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=97830 $D=1
M403 437 73 237 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=102460 $D=1
M404 5 436 750 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=97830 $D=1
M405 5 437 751 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=102460 $D=1
M406 438 750 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=97830 $D=1
M407 439 751 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=102460 $D=1
M408 436 432 438 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=97830 $D=1
M409 437 433 439 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=102460 $D=1
M410 438 74 246 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=97830 $D=1
M411 439 74 247 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=102460 $D=1
M412 250 75 438 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=97830 $D=1
M413 251 75 439 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=102460 $D=1
M414 440 75 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=97830 $D=1
M415 441 75 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=102460 $D=1
M416 5 76 442 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=97830 $D=1
M417 5 76 443 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=102460 $D=1
M418 444 77 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=97830 $D=1
M419 445 77 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=102460 $D=1
M420 446 76 236 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=97830 $D=1
M421 447 76 237 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=102460 $D=1
M422 5 446 752 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=97830 $D=1
M423 5 447 753 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=102460 $D=1
M424 448 752 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=97830 $D=1
M425 449 753 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=102460 $D=1
M426 446 442 448 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=97830 $D=1
M427 447 443 449 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=102460 $D=1
M428 448 77 246 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=97830 $D=1
M429 449 77 247 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=102460 $D=1
M430 250 78 448 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=97830 $D=1
M431 251 78 449 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=102460 $D=1
M432 450 78 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=97830 $D=1
M433 451 78 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=102460 $D=1
M434 5 79 452 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=97830 $D=1
M435 5 79 453 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=102460 $D=1
M436 454 80 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=97830 $D=1
M437 455 80 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=102460 $D=1
M438 456 79 236 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=97830 $D=1
M439 457 79 237 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=102460 $D=1
M440 5 456 754 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=97830 $D=1
M441 5 457 755 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=102460 $D=1
M442 458 754 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=97830 $D=1
M443 459 755 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=102460 $D=1
M444 456 452 458 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=97830 $D=1
M445 457 453 459 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=102460 $D=1
M446 458 80 246 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=97830 $D=1
M447 459 80 247 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=102460 $D=1
M448 250 81 458 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=97830 $D=1
M449 251 81 459 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=102460 $D=1
M450 460 81 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=97830 $D=1
M451 461 81 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=102460 $D=1
M452 5 82 462 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=97830 $D=1
M453 5 82 463 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=102460 $D=1
M454 464 83 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=97830 $D=1
M455 465 83 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=102460 $D=1
M456 466 82 236 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=97830 $D=1
M457 467 82 237 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=102460 $D=1
M458 5 466 756 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=97830 $D=1
M459 5 467 757 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=102460 $D=1
M460 468 756 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=97830 $D=1
M461 469 757 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=102460 $D=1
M462 466 462 468 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=97830 $D=1
M463 467 463 469 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=102460 $D=1
M464 468 83 246 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=97830 $D=1
M465 469 83 247 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=102460 $D=1
M466 250 84 468 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=97830 $D=1
M467 251 84 469 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=102460 $D=1
M468 470 84 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=97830 $D=1
M469 471 84 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=102460 $D=1
M470 5 85 472 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=97830 $D=1
M471 5 85 473 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=102460 $D=1
M472 474 86 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=97830 $D=1
M473 475 86 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=102460 $D=1
M474 476 85 236 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=97830 $D=1
M475 477 85 237 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=102460 $D=1
M476 5 476 758 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=97830 $D=1
M477 5 477 759 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=102460 $D=1
M478 478 758 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=97830 $D=1
M479 479 759 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=102460 $D=1
M480 476 472 478 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=97830 $D=1
M481 477 473 479 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=102460 $D=1
M482 478 86 246 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=97830 $D=1
M483 479 86 247 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=102460 $D=1
M484 250 87 478 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=97830 $D=1
M485 251 87 479 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=102460 $D=1
M486 480 87 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=97830 $D=1
M487 481 87 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=102460 $D=1
M488 5 88 482 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=97830 $D=1
M489 5 88 483 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=102460 $D=1
M490 484 89 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=97830 $D=1
M491 485 89 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=102460 $D=1
M492 486 88 236 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=97830 $D=1
M493 487 88 237 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=102460 $D=1
M494 5 486 760 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=97830 $D=1
M495 5 487 761 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=102460 $D=1
M496 488 760 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=97830 $D=1
M497 489 761 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=102460 $D=1
M498 486 482 488 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=97830 $D=1
M499 487 483 489 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=102460 $D=1
M500 488 89 246 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=97830 $D=1
M501 489 89 247 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=102460 $D=1
M502 250 90 488 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=97830 $D=1
M503 251 90 489 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=102460 $D=1
M504 490 90 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=97830 $D=1
M505 491 90 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=102460 $D=1
M506 5 91 492 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=97830 $D=1
M507 5 91 493 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=102460 $D=1
M508 494 92 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=97830 $D=1
M509 495 92 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=102460 $D=1
M510 496 91 236 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=97830 $D=1
M511 497 91 237 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=102460 $D=1
M512 5 496 762 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=97830 $D=1
M513 5 497 763 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=102460 $D=1
M514 498 762 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=97830 $D=1
M515 499 763 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=102460 $D=1
M516 496 492 498 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=97830 $D=1
M517 497 493 499 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=102460 $D=1
M518 498 92 246 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=97830 $D=1
M519 499 92 247 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=102460 $D=1
M520 250 93 498 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=97830 $D=1
M521 251 93 499 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=102460 $D=1
M522 500 93 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=97830 $D=1
M523 501 93 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=102460 $D=1
M524 5 94 502 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=97830 $D=1
M525 5 94 503 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=102460 $D=1
M526 504 95 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=97830 $D=1
M527 505 95 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=102460 $D=1
M528 506 94 236 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=97830 $D=1
M529 507 94 237 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=102460 $D=1
M530 5 506 764 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=97830 $D=1
M531 5 507 765 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=102460 $D=1
M532 508 764 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=97830 $D=1
M533 509 765 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=102460 $D=1
M534 506 502 508 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=97830 $D=1
M535 507 503 509 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=102460 $D=1
M536 508 95 246 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=97830 $D=1
M537 509 95 247 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=102460 $D=1
M538 250 96 508 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=97830 $D=1
M539 251 96 509 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=102460 $D=1
M540 510 96 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=97830 $D=1
M541 511 96 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=102460 $D=1
M542 5 97 512 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=97830 $D=1
M543 5 97 513 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=102460 $D=1
M544 514 98 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=97830 $D=1
M545 515 98 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=102460 $D=1
M546 516 97 236 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=97830 $D=1
M547 517 97 237 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=102460 $D=1
M548 5 516 766 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=97830 $D=1
M549 5 517 767 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=102460 $D=1
M550 518 766 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=97830 $D=1
M551 519 767 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=102460 $D=1
M552 516 512 518 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=97830 $D=1
M553 517 513 519 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=102460 $D=1
M554 518 98 246 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=97830 $D=1
M555 519 98 247 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=102460 $D=1
M556 250 99 518 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=97830 $D=1
M557 251 99 519 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=102460 $D=1
M558 520 99 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=97830 $D=1
M559 521 99 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=102460 $D=1
M560 5 100 522 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=97830 $D=1
M561 5 100 523 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=102460 $D=1
M562 524 101 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=97830 $D=1
M563 525 101 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=102460 $D=1
M564 526 100 236 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=97830 $D=1
M565 527 100 237 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=102460 $D=1
M566 5 526 768 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=97830 $D=1
M567 5 527 769 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=102460 $D=1
M568 528 768 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=97830 $D=1
M569 529 769 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=102460 $D=1
M570 526 522 528 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=97830 $D=1
M571 527 523 529 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=102460 $D=1
M572 528 101 246 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=97830 $D=1
M573 529 101 247 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=102460 $D=1
M574 250 102 528 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=97830 $D=1
M575 251 102 529 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=102460 $D=1
M576 530 102 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=97830 $D=1
M577 531 102 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=102460 $D=1
M578 5 103 532 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=97830 $D=1
M579 5 103 533 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=102460 $D=1
M580 534 104 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=97830 $D=1
M581 535 104 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=102460 $D=1
M582 536 103 236 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=97830 $D=1
M583 537 103 237 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=102460 $D=1
M584 5 536 770 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=97830 $D=1
M585 5 537 771 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=102460 $D=1
M586 538 770 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=97830 $D=1
M587 539 771 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=102460 $D=1
M588 536 532 538 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=97830 $D=1
M589 537 533 539 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=102460 $D=1
M590 538 104 246 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=97830 $D=1
M591 539 104 247 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=102460 $D=1
M592 250 105 538 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=97830 $D=1
M593 251 105 539 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=102460 $D=1
M594 540 105 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=97830 $D=1
M595 541 105 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=102460 $D=1
M596 5 106 542 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=97830 $D=1
M597 5 106 543 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=102460 $D=1
M598 544 107 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=97830 $D=1
M599 545 107 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=102460 $D=1
M600 546 106 236 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=97830 $D=1
M601 547 106 237 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=102460 $D=1
M602 5 546 772 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=97830 $D=1
M603 5 547 773 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=102460 $D=1
M604 548 772 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=97830 $D=1
M605 549 773 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=102460 $D=1
M606 546 542 548 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=97830 $D=1
M607 547 543 549 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=102460 $D=1
M608 548 107 246 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=97830 $D=1
M609 549 107 247 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=102460 $D=1
M610 250 108 548 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=97830 $D=1
M611 251 108 549 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=102460 $D=1
M612 550 108 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=97830 $D=1
M613 551 108 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=102460 $D=1
M614 5 109 552 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=97830 $D=1
M615 5 109 553 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=102460 $D=1
M616 554 110 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=97830 $D=1
M617 555 110 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=102460 $D=1
M618 5 110 246 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=97830 $D=1
M619 5 110 247 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=102460 $D=1
M620 250 109 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=97830 $D=1
M621 251 109 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=102460 $D=1
M622 5 558 556 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=97830 $D=1
M623 5 559 557 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=102460 $D=1
M624 558 111 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=97830 $D=1
M625 559 111 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=102460 $D=1
M626 774 246 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=97830 $D=1
M627 775 247 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=102460 $D=1
M628 560 556 774 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=97830 $D=1
M629 561 557 775 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=102460 $D=1
M630 5 560 562 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=97830 $D=1
M631 5 561 563 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=102460 $D=1
M632 776 562 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=97830 $D=1
M633 777 563 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=102460 $D=1
M634 560 558 776 5 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=97830 $D=1
M635 561 559 777 5 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=102460 $D=1
M636 5 566 564 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=97830 $D=1
M637 5 567 565 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=102460 $D=1
M638 566 111 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=97830 $D=1
M639 567 111 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=102460 $D=1
M640 778 250 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=97830 $D=1
M641 779 251 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=102460 $D=1
M642 568 564 778 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=97830 $D=1
M643 569 565 779 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=102460 $D=1
M644 5 568 112 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=97830 $D=1
M645 5 569 113 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=102460 $D=1
M646 780 112 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=97830 $D=1
M647 781 113 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=102460 $D=1
M648 568 566 780 5 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=97830 $D=1
M649 569 567 781 5 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=102460 $D=1
M650 570 115 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=97830 $D=1
M651 571 115 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=102460 $D=1
M652 572 570 562 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=97830 $D=1
M653 573 571 563 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=102460 $D=1
M654 117 115 572 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=97830 $D=1
M655 118 115 573 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=102460 $D=1
M656 574 119 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=97830 $D=1
M657 575 119 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=102460 $D=1
M658 576 574 112 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=97830 $D=1
M659 577 575 113 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=102460 $D=1
M660 782 119 576 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=97830 $D=1
M661 783 119 577 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=102460 $D=1
M662 5 112 782 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=97830 $D=1
M663 5 113 783 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=102460 $D=1
M664 578 122 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=97830 $D=1
M665 579 122 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=102460 $D=1
M666 580 578 576 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=97830 $D=1
M667 581 579 577 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=102460 $D=1
M668 10 122 580 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=97830 $D=1
M669 11 122 581 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=102460 $D=1
M670 583 582 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=97830 $D=1
M671 584 123 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=102460 $D=1
M672 5 587 585 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=97830 $D=1
M673 5 588 586 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=102460 $D=1
M674 589 572 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=97830 $D=1
M675 590 573 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=102460 $D=1
M676 587 589 582 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=97830 $D=1
M677 588 590 123 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=102460 $D=1
M678 583 572 587 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=97830 $D=1
M679 584 573 588 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=102460 $D=1
M680 591 585 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=97830 $D=1
M681 592 586 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=102460 $D=1
M682 126 591 580 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=97830 $D=1
M683 582 592 581 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=102460 $D=1
M684 572 585 126 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=97830 $D=1
M685 573 586 582 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=102460 $D=1
M686 593 126 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=97830 $D=1
M687 594 582 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=102460 $D=1
M688 595 585 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=97830 $D=1
M689 596 586 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=102460 $D=1
M690 597 595 593 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=97830 $D=1
M691 598 596 594 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=102460 $D=1
M692 580 585 597 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=97830 $D=1
M693 581 586 598 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=102460 $D=1
M694 599 572 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=97830 $D=1
M695 600 573 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=102460 $D=1
M696 5 580 599 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=97830 $D=1
M697 5 581 600 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=102460 $D=1
M698 601 597 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=97830 $D=1
M699 602 598 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=102460 $D=1
M700 802 572 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=97830 $D=1
M701 803 573 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=102460 $D=1
M702 603 580 802 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=97830 $D=1
M703 604 581 803 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=102460 $D=1
M704 804 572 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=97830 $D=1
M705 805 573 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=102460 $D=1
M706 605 580 804 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=97830 $D=1
M707 606 581 805 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=102460 $D=1
M708 609 572 607 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=97830 $D=1
M709 610 573 608 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=102460 $D=1
M710 607 580 609 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=97830 $D=1
M711 608 581 610 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=102460 $D=1
M712 5 605 607 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=97830 $D=1
M713 5 606 608 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=102460 $D=1
M714 611 128 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=97830 $D=1
M715 612 128 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=102460 $D=1
M716 613 611 599 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=97830 $D=1
M717 614 612 600 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=102460 $D=1
M718 603 128 613 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=97830 $D=1
M719 604 128 614 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=102460 $D=1
M720 615 611 601 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=97830 $D=1
M721 616 612 602 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=102460 $D=1
M722 609 128 615 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=97830 $D=1
M723 610 128 616 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=102460 $D=1
M724 617 129 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=97830 $D=1
M725 618 129 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=102460 $D=1
M726 619 617 615 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=97830 $D=1
M727 620 618 616 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=102460 $D=1
M728 613 129 619 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=97830 $D=1
M729 614 129 620 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=102460 $D=1
M730 12 619 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=97830 $D=1
M731 13 620 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=102460 $D=1
M732 621 130 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=97830 $D=1
M733 622 130 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=102460 $D=1
M734 623 621 131 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=97830 $D=1
M735 624 622 132 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=102460 $D=1
M736 133 130 623 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=97830 $D=1
M737 134 130 624 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=102460 $D=1
M738 625 130 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=97830 $D=1
M739 626 130 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=102460 $D=1
M740 627 625 135 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=97830 $D=1
M741 628 626 136 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=102460 $D=1
M742 137 130 627 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=97830 $D=1
M743 138 130 628 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=102460 $D=1
M744 629 130 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=97830 $D=1
M745 630 130 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=102460 $D=1
M746 631 629 139 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=97830 $D=1
M747 632 630 140 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=102460 $D=1
M748 116 130 631 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=97830 $D=1
M749 121 130 632 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=102460 $D=1
M750 633 130 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=97830 $D=1
M751 634 130 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=102460 $D=1
M752 635 633 141 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=97830 $D=1
M753 636 634 142 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=102460 $D=1
M754 114 130 635 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=97830 $D=1
M755 120 130 636 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=102460 $D=1
M756 637 130 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=97830 $D=1
M757 638 130 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=102460 $D=1
M758 639 637 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=97830 $D=1
M759 640 638 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=102460 $D=1
M760 143 130 639 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=97830 $D=1
M761 144 130 640 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=102460 $D=1
M762 5 572 784 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=97830 $D=1
M763 5 573 785 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=102460 $D=1
M764 134 784 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=97830 $D=1
M765 131 785 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=102460 $D=1
M766 641 145 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=97830 $D=1
M767 642 145 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=102460 $D=1
M768 146 641 134 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=97830 $D=1
M769 147 642 131 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=102460 $D=1
M770 623 145 146 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=97830 $D=1
M771 624 145 147 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=102460 $D=1
M772 643 148 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=97830 $D=1
M773 644 148 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=102460 $D=1
M774 149 643 146 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=97830 $D=1
M775 127 644 147 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=102460 $D=1
M776 627 148 149 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=97830 $D=1
M777 628 148 127 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=102460 $D=1
M778 645 150 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=97830 $D=1
M779 646 150 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=102460 $D=1
M780 124 645 149 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=97830 $D=1
M781 125 646 127 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=102460 $D=1
M782 631 150 124 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=97830 $D=1
M783 632 150 125 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=102460 $D=1
M784 647 151 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=97830 $D=1
M785 648 151 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=102460 $D=1
M786 152 647 124 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=97830 $D=1
M787 153 648 125 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=102460 $D=1
M788 635 151 152 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=97830 $D=1
M789 636 151 153 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=102460 $D=1
M790 649 154 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=97830 $D=1
M791 650 154 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=102460 $D=1
M792 222 649 152 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=97830 $D=1
M793 223 650 153 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=102460 $D=1
M794 639 154 222 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=97830 $D=1
M795 640 154 223 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=102460 $D=1
M796 651 155 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=97830 $D=1
M797 652 155 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=102460 $D=1
M798 653 651 112 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=97830 $D=1
M799 654 652 113 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=102460 $D=1
M800 10 155 653 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=97830 $D=1
M801 11 155 654 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=102460 $D=1
M802 806 562 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=97830 $D=1
M803 807 563 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=102460 $D=1
M804 655 653 806 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=97830 $D=1
M805 656 654 807 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=102460 $D=1
M806 659 562 657 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=97830 $D=1
M807 660 563 658 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=102460 $D=1
M808 657 653 659 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=97830 $D=1
M809 658 654 660 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=102460 $D=1
M810 5 655 657 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=97830 $D=1
M811 5 656 658 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=102460 $D=1
M812 808 156 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=97830 $D=1
M813 809 661 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=102460 $D=1
M814 786 659 808 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=97830 $D=1
M815 787 660 809 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=102460 $D=1
M816 661 786 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=97830 $D=1
M817 157 787 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=102460 $D=1
M818 662 562 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=97830 $D=1
M819 663 563 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=102460 $D=1
M820 5 664 662 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=97830 $D=1
M821 5 665 663 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=102460 $D=1
M822 664 653 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=97830 $D=1
M823 665 654 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=102460 $D=1
M824 810 662 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=97830 $D=1
M825 811 663 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=102460 $D=1
M826 666 156 810 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=97830 $D=1
M827 667 661 811 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=102460 $D=1
M828 669 158 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=97830 $D=1
M829 670 668 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=102460 $D=1
M830 812 666 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=97830 $D=1
M831 813 667 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=102460 $D=1
M832 668 669 812 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=97830 $D=1
M833 159 670 813 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=102460 $D=1
M834 672 671 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=97830 $D=1
M835 673 160 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=102460 $D=1
M836 5 676 674 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=97830 $D=1
M837 5 677 675 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=102460 $D=1
M838 678 117 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=97830 $D=1
M839 679 118 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=102460 $D=1
M840 676 678 671 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=97830 $D=1
M841 677 679 160 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=102460 $D=1
M842 672 117 676 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=97830 $D=1
M843 673 118 677 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=102460 $D=1
M844 680 674 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=97830 $D=1
M845 681 675 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=102460 $D=1
M846 161 680 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=97830 $D=1
M847 671 681 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=102460 $D=1
M848 117 674 161 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=97830 $D=1
M849 118 675 671 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=102460 $D=1
M850 682 161 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=97830 $D=1
M851 683 671 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=102460 $D=1
M852 684 674 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=97830 $D=1
M853 685 675 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=102460 $D=1
M854 224 684 682 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=97830 $D=1
M855 225 685 683 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=102460 $D=1
M856 5 674 224 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=97830 $D=1
M857 5 675 225 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=102460 $D=1
M858 686 162 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=97830 $D=1
M859 687 162 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=102460 $D=1
M860 688 686 224 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=97830 $D=1
M861 689 687 225 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=102460 $D=1
M862 12 162 688 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=97830 $D=1
M863 13 162 689 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=102460 $D=1
M864 690 163 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=97830 $D=1
M865 691 163 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=102460 $D=1
M866 692 690 688 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=97830 $D=1
M867 693 691 689 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=102460 $D=1
M868 5 163 692 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=97830 $D=1
M869 5 163 693 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=102460 $D=1
M870 694 111 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=97830 $D=1
M871 695 111 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=102460 $D=1
M872 5 694 696 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=97830 $D=1
M873 5 695 697 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=102460 $D=1
M874 698 111 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=97830 $D=1
M875 699 111 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=102460 $D=1
M876 700 694 692 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=97830 $D=1
M877 701 695 693 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=102460 $D=1
M878 5 700 788 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=97830 $D=1
M879 5 701 789 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=102460 $D=1
M880 702 788 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=97830 $D=1
M881 703 789 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=102460 $D=1
M882 700 696 702 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=97830 $D=1
M883 701 697 703 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=102460 $D=1
M884 704 111 702 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=97830 $D=1
M885 705 111 703 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=102460 $D=1
M886 5 708 706 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=97830 $D=1
M887 5 709 707 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=102460 $D=1
M888 708 111 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=97830 $D=1
M889 709 111 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=102460 $D=1
M890 790 704 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=97830 $D=1
M891 791 705 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=102460 $D=1
M892 710 706 790 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=97830 $D=1
M893 711 707 791 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=102460 $D=1
M894 5 710 117 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=97830 $D=1
M895 5 711 118 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=102460 $D=1
M896 792 117 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=97830 $D=1
M897 793 118 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=102460 $D=1
M898 710 708 792 5 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=97830 $D=1
M899 711 709 793 5 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=102460 $D=1
M900 198 1 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=99080 $D=0
M901 199 1 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=103710 $D=0
M902 200 1 2 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=99080 $D=0
M903 201 1 3 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=103710 $D=0
M904 5 198 200 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=99080 $D=0
M905 5 199 201 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=103710 $D=0
M906 202 1 4 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=99080 $D=0
M907 203 1 4 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=103710 $D=0
M908 2 198 202 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=99080 $D=0
M909 3 199 203 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=103710 $D=0
M910 204 1 5 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=99080 $D=0
M911 205 1 5 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=103710 $D=0
M912 2 198 204 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=99080 $D=0
M913 3 199 205 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=103710 $D=0
M914 208 6 204 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=99080 $D=0
M915 209 6 205 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=103710 $D=0
M916 206 6 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=99080 $D=0
M917 207 6 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=103710 $D=0
M918 210 6 202 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=99080 $D=0
M919 211 6 203 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=103710 $D=0
M920 200 206 210 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=99080 $D=0
M921 201 207 211 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=103710 $D=0
M922 212 7 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=99080 $D=0
M923 213 7 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=103710 $D=0
M924 214 7 210 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=99080 $D=0
M925 215 7 211 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=103710 $D=0
M926 208 212 214 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=99080 $D=0
M927 209 213 215 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=103710 $D=0
M928 216 9 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=99080 $D=0
M929 217 9 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=103710 $D=0
M930 218 9 5 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=99080 $D=0
M931 219 9 5 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=103710 $D=0
M932 10 216 218 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=99080 $D=0
M933 11 217 219 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=103710 $D=0
M934 220 9 12 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=99080 $D=0
M935 221 9 13 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=103710 $D=0
M936 222 216 220 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=99080 $D=0
M937 223 217 221 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=103710 $D=0
M938 226 9 224 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=99080 $D=0
M939 227 9 225 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=103710 $D=0
M940 214 216 226 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=99080 $D=0
M941 215 217 227 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=103710 $D=0
M942 230 14 226 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=99080 $D=0
M943 231 14 227 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=103710 $D=0
M944 228 14 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=99080 $D=0
M945 229 14 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=103710 $D=0
M946 232 14 220 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=99080 $D=0
M947 233 14 221 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=103710 $D=0
M948 218 228 232 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=99080 $D=0
M949 219 229 233 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=103710 $D=0
M950 234 15 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=99080 $D=0
M951 235 15 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=103710 $D=0
M952 236 15 232 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=99080 $D=0
M953 237 15 233 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=103710 $D=0
M954 230 234 236 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=99080 $D=0
M955 231 235 237 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=103710 $D=0
M956 8 16 238 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=99080 $D=0
M957 8 16 239 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=103710 $D=0
M958 240 17 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=99080 $D=0
M959 241 17 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=103710 $D=0
M960 242 238 236 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=99080 $D=0
M961 243 239 237 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=103710 $D=0
M962 8 242 712 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=99080 $D=0
M963 8 243 713 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=103710 $D=0
M964 244 712 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=99080 $D=0
M965 245 713 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=103710 $D=0
M966 242 16 244 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=99080 $D=0
M967 243 16 245 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=103710 $D=0
M968 244 240 246 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=99080 $D=0
M969 245 241 247 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=103710 $D=0
M970 250 248 244 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=99080 $D=0
M971 251 249 245 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=103710 $D=0
M972 248 18 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=99080 $D=0
M973 249 18 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=103710 $D=0
M974 8 19 252 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=99080 $D=0
M975 8 19 253 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=103710 $D=0
M976 254 20 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=99080 $D=0
M977 255 20 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=103710 $D=0
M978 256 252 236 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=99080 $D=0
M979 257 253 237 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=103710 $D=0
M980 8 256 714 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=99080 $D=0
M981 8 257 715 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=103710 $D=0
M982 258 714 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=99080 $D=0
M983 259 715 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=103710 $D=0
M984 256 19 258 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=99080 $D=0
M985 257 19 259 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=103710 $D=0
M986 258 254 246 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=99080 $D=0
M987 259 255 247 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=103710 $D=0
M988 250 260 258 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=99080 $D=0
M989 251 261 259 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=103710 $D=0
M990 260 21 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=99080 $D=0
M991 261 21 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=103710 $D=0
M992 8 22 262 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=99080 $D=0
M993 8 22 263 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=103710 $D=0
M994 264 23 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=99080 $D=0
M995 265 23 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=103710 $D=0
M996 266 262 236 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=99080 $D=0
M997 267 263 237 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=103710 $D=0
M998 8 266 716 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=99080 $D=0
M999 8 267 717 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=103710 $D=0
M1000 268 716 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=99080 $D=0
M1001 269 717 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=103710 $D=0
M1002 266 22 268 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=99080 $D=0
M1003 267 22 269 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=103710 $D=0
M1004 268 264 246 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=99080 $D=0
M1005 269 265 247 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=103710 $D=0
M1006 250 270 268 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=99080 $D=0
M1007 251 271 269 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=103710 $D=0
M1008 270 24 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=99080 $D=0
M1009 271 24 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=103710 $D=0
M1010 8 25 272 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=99080 $D=0
M1011 8 25 273 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=103710 $D=0
M1012 274 26 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=99080 $D=0
M1013 275 26 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=103710 $D=0
M1014 276 272 236 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=99080 $D=0
M1015 277 273 237 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=103710 $D=0
M1016 8 276 718 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=99080 $D=0
M1017 8 277 719 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=103710 $D=0
M1018 278 718 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=99080 $D=0
M1019 279 719 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=103710 $D=0
M1020 276 25 278 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=99080 $D=0
M1021 277 25 279 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=103710 $D=0
M1022 278 274 246 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=99080 $D=0
M1023 279 275 247 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=103710 $D=0
M1024 250 280 278 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=99080 $D=0
M1025 251 281 279 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=103710 $D=0
M1026 280 27 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=99080 $D=0
M1027 281 27 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=103710 $D=0
M1028 8 28 282 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=99080 $D=0
M1029 8 28 283 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=103710 $D=0
M1030 284 29 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=99080 $D=0
M1031 285 29 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=103710 $D=0
M1032 286 282 236 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=99080 $D=0
M1033 287 283 237 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=103710 $D=0
M1034 8 286 720 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=99080 $D=0
M1035 8 287 721 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=103710 $D=0
M1036 288 720 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=99080 $D=0
M1037 289 721 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=103710 $D=0
M1038 286 28 288 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=99080 $D=0
M1039 287 28 289 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=103710 $D=0
M1040 288 284 246 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=99080 $D=0
M1041 289 285 247 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=103710 $D=0
M1042 250 290 288 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=99080 $D=0
M1043 251 291 289 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=103710 $D=0
M1044 290 30 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=99080 $D=0
M1045 291 30 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=103710 $D=0
M1046 8 31 292 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=99080 $D=0
M1047 8 31 293 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=103710 $D=0
M1048 294 32 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=99080 $D=0
M1049 295 32 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=103710 $D=0
M1050 296 292 236 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=99080 $D=0
M1051 297 293 237 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=103710 $D=0
M1052 8 296 722 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=99080 $D=0
M1053 8 297 723 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=103710 $D=0
M1054 298 722 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=99080 $D=0
M1055 299 723 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=103710 $D=0
M1056 296 31 298 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=99080 $D=0
M1057 297 31 299 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=103710 $D=0
M1058 298 294 246 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=99080 $D=0
M1059 299 295 247 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=103710 $D=0
M1060 250 300 298 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=99080 $D=0
M1061 251 301 299 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=103710 $D=0
M1062 300 33 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=99080 $D=0
M1063 301 33 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=103710 $D=0
M1064 8 34 302 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=99080 $D=0
M1065 8 34 303 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=103710 $D=0
M1066 304 35 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=99080 $D=0
M1067 305 35 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=103710 $D=0
M1068 306 302 236 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=99080 $D=0
M1069 307 303 237 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=103710 $D=0
M1070 8 306 724 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=99080 $D=0
M1071 8 307 725 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=103710 $D=0
M1072 308 724 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=99080 $D=0
M1073 309 725 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=103710 $D=0
M1074 306 34 308 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=99080 $D=0
M1075 307 34 309 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=103710 $D=0
M1076 308 304 246 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=99080 $D=0
M1077 309 305 247 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=103710 $D=0
M1078 250 310 308 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=99080 $D=0
M1079 251 311 309 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=103710 $D=0
M1080 310 36 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=99080 $D=0
M1081 311 36 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=103710 $D=0
M1082 8 37 312 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=99080 $D=0
M1083 8 37 313 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=103710 $D=0
M1084 314 38 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=99080 $D=0
M1085 315 38 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=103710 $D=0
M1086 316 312 236 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=99080 $D=0
M1087 317 313 237 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=103710 $D=0
M1088 8 316 726 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=99080 $D=0
M1089 8 317 727 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=103710 $D=0
M1090 318 726 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=99080 $D=0
M1091 319 727 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=103710 $D=0
M1092 316 37 318 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=99080 $D=0
M1093 317 37 319 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=103710 $D=0
M1094 318 314 246 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=99080 $D=0
M1095 319 315 247 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=103710 $D=0
M1096 250 320 318 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=99080 $D=0
M1097 251 321 319 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=103710 $D=0
M1098 320 39 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=99080 $D=0
M1099 321 39 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=103710 $D=0
M1100 8 40 322 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=99080 $D=0
M1101 8 40 323 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=103710 $D=0
M1102 324 41 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=99080 $D=0
M1103 325 41 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=103710 $D=0
M1104 326 322 236 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=99080 $D=0
M1105 327 323 237 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=103710 $D=0
M1106 8 326 728 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=99080 $D=0
M1107 8 327 729 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=103710 $D=0
M1108 328 728 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=99080 $D=0
M1109 329 729 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=103710 $D=0
M1110 326 40 328 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=99080 $D=0
M1111 327 40 329 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=103710 $D=0
M1112 328 324 246 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=99080 $D=0
M1113 329 325 247 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=103710 $D=0
M1114 250 330 328 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=99080 $D=0
M1115 251 331 329 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=103710 $D=0
M1116 330 42 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=99080 $D=0
M1117 331 42 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=103710 $D=0
M1118 8 43 332 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=99080 $D=0
M1119 8 43 333 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=103710 $D=0
M1120 334 44 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=99080 $D=0
M1121 335 44 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=103710 $D=0
M1122 336 332 236 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=99080 $D=0
M1123 337 333 237 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=103710 $D=0
M1124 8 336 730 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=99080 $D=0
M1125 8 337 731 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=103710 $D=0
M1126 338 730 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=99080 $D=0
M1127 339 731 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=103710 $D=0
M1128 336 43 338 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=99080 $D=0
M1129 337 43 339 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=103710 $D=0
M1130 338 334 246 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=99080 $D=0
M1131 339 335 247 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=103710 $D=0
M1132 250 340 338 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=99080 $D=0
M1133 251 341 339 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=103710 $D=0
M1134 340 45 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=99080 $D=0
M1135 341 45 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=103710 $D=0
M1136 8 46 342 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=99080 $D=0
M1137 8 46 343 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=103710 $D=0
M1138 344 47 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=99080 $D=0
M1139 345 47 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=103710 $D=0
M1140 346 342 236 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=99080 $D=0
M1141 347 343 237 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=103710 $D=0
M1142 8 346 732 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=99080 $D=0
M1143 8 347 733 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=103710 $D=0
M1144 348 732 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=99080 $D=0
M1145 349 733 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=103710 $D=0
M1146 346 46 348 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=99080 $D=0
M1147 347 46 349 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=103710 $D=0
M1148 348 344 246 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=99080 $D=0
M1149 349 345 247 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=103710 $D=0
M1150 250 350 348 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=99080 $D=0
M1151 251 351 349 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=103710 $D=0
M1152 350 48 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=99080 $D=0
M1153 351 48 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=103710 $D=0
M1154 8 49 352 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=99080 $D=0
M1155 8 49 353 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=103710 $D=0
M1156 354 50 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=99080 $D=0
M1157 355 50 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=103710 $D=0
M1158 356 352 236 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=99080 $D=0
M1159 357 353 237 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=103710 $D=0
M1160 8 356 734 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=99080 $D=0
M1161 8 357 735 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=103710 $D=0
M1162 358 734 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=99080 $D=0
M1163 359 735 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=103710 $D=0
M1164 356 49 358 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=99080 $D=0
M1165 357 49 359 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=103710 $D=0
M1166 358 354 246 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=99080 $D=0
M1167 359 355 247 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=103710 $D=0
M1168 250 360 358 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=99080 $D=0
M1169 251 361 359 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=103710 $D=0
M1170 360 51 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=99080 $D=0
M1171 361 51 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=103710 $D=0
M1172 8 52 362 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=99080 $D=0
M1173 8 52 363 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=103710 $D=0
M1174 364 53 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=99080 $D=0
M1175 365 53 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=103710 $D=0
M1176 366 362 236 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=99080 $D=0
M1177 367 363 237 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=103710 $D=0
M1178 8 366 736 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=99080 $D=0
M1179 8 367 737 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=103710 $D=0
M1180 368 736 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=99080 $D=0
M1181 369 737 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=103710 $D=0
M1182 366 52 368 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=99080 $D=0
M1183 367 52 369 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=103710 $D=0
M1184 368 364 246 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=99080 $D=0
M1185 369 365 247 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=103710 $D=0
M1186 250 370 368 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=99080 $D=0
M1187 251 371 369 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=103710 $D=0
M1188 370 54 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=99080 $D=0
M1189 371 54 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=103710 $D=0
M1190 8 55 372 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=99080 $D=0
M1191 8 55 373 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=103710 $D=0
M1192 374 56 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=99080 $D=0
M1193 375 56 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=103710 $D=0
M1194 376 372 236 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=99080 $D=0
M1195 377 373 237 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=103710 $D=0
M1196 8 376 738 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=99080 $D=0
M1197 8 377 739 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=103710 $D=0
M1198 378 738 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=99080 $D=0
M1199 379 739 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=103710 $D=0
M1200 376 55 378 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=99080 $D=0
M1201 377 55 379 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=103710 $D=0
M1202 378 374 246 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=99080 $D=0
M1203 379 375 247 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=103710 $D=0
M1204 250 380 378 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=99080 $D=0
M1205 251 381 379 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=103710 $D=0
M1206 380 57 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=99080 $D=0
M1207 381 57 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=103710 $D=0
M1208 8 58 382 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=99080 $D=0
M1209 8 58 383 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=103710 $D=0
M1210 384 59 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=99080 $D=0
M1211 385 59 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=103710 $D=0
M1212 386 382 236 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=99080 $D=0
M1213 387 383 237 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=103710 $D=0
M1214 8 386 740 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=99080 $D=0
M1215 8 387 741 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=103710 $D=0
M1216 388 740 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=99080 $D=0
M1217 389 741 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=103710 $D=0
M1218 386 58 388 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=99080 $D=0
M1219 387 58 389 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=103710 $D=0
M1220 388 384 246 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=99080 $D=0
M1221 389 385 247 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=103710 $D=0
M1222 250 390 388 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=99080 $D=0
M1223 251 391 389 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=103710 $D=0
M1224 390 60 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=99080 $D=0
M1225 391 60 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=103710 $D=0
M1226 8 61 392 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=99080 $D=0
M1227 8 61 393 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=103710 $D=0
M1228 394 62 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=99080 $D=0
M1229 395 62 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=103710 $D=0
M1230 396 392 236 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=99080 $D=0
M1231 397 393 237 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=103710 $D=0
M1232 8 396 742 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=99080 $D=0
M1233 8 397 743 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=103710 $D=0
M1234 398 742 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=99080 $D=0
M1235 399 743 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=103710 $D=0
M1236 396 61 398 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=99080 $D=0
M1237 397 61 399 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=103710 $D=0
M1238 398 394 246 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=99080 $D=0
M1239 399 395 247 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=103710 $D=0
M1240 250 400 398 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=99080 $D=0
M1241 251 401 399 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=103710 $D=0
M1242 400 63 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=99080 $D=0
M1243 401 63 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=103710 $D=0
M1244 8 64 402 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=99080 $D=0
M1245 8 64 403 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=103710 $D=0
M1246 404 65 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=99080 $D=0
M1247 405 65 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=103710 $D=0
M1248 406 402 236 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=99080 $D=0
M1249 407 403 237 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=103710 $D=0
M1250 8 406 744 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=99080 $D=0
M1251 8 407 745 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=103710 $D=0
M1252 408 744 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=99080 $D=0
M1253 409 745 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=103710 $D=0
M1254 406 64 408 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=99080 $D=0
M1255 407 64 409 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=103710 $D=0
M1256 408 404 246 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=99080 $D=0
M1257 409 405 247 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=103710 $D=0
M1258 250 410 408 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=99080 $D=0
M1259 251 411 409 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=103710 $D=0
M1260 410 66 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=99080 $D=0
M1261 411 66 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=103710 $D=0
M1262 8 67 412 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=99080 $D=0
M1263 8 67 413 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=103710 $D=0
M1264 414 68 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=99080 $D=0
M1265 415 68 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=103710 $D=0
M1266 416 412 236 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=99080 $D=0
M1267 417 413 237 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=103710 $D=0
M1268 8 416 746 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=99080 $D=0
M1269 8 417 747 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=103710 $D=0
M1270 418 746 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=99080 $D=0
M1271 419 747 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=103710 $D=0
M1272 416 67 418 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=99080 $D=0
M1273 417 67 419 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=103710 $D=0
M1274 418 414 246 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=99080 $D=0
M1275 419 415 247 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=103710 $D=0
M1276 250 420 418 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=99080 $D=0
M1277 251 421 419 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=103710 $D=0
M1278 420 69 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=99080 $D=0
M1279 421 69 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=103710 $D=0
M1280 8 70 422 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=99080 $D=0
M1281 8 70 423 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=103710 $D=0
M1282 424 71 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=99080 $D=0
M1283 425 71 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=103710 $D=0
M1284 426 422 236 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=99080 $D=0
M1285 427 423 237 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=103710 $D=0
M1286 8 426 748 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=99080 $D=0
M1287 8 427 749 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=103710 $D=0
M1288 428 748 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=99080 $D=0
M1289 429 749 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=103710 $D=0
M1290 426 70 428 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=99080 $D=0
M1291 427 70 429 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=103710 $D=0
M1292 428 424 246 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=99080 $D=0
M1293 429 425 247 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=103710 $D=0
M1294 250 430 428 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=99080 $D=0
M1295 251 431 429 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=103710 $D=0
M1296 430 72 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=99080 $D=0
M1297 431 72 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=103710 $D=0
M1298 8 73 432 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=99080 $D=0
M1299 8 73 433 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=103710 $D=0
M1300 434 74 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=99080 $D=0
M1301 435 74 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=103710 $D=0
M1302 436 432 236 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=99080 $D=0
M1303 437 433 237 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=103710 $D=0
M1304 8 436 750 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=99080 $D=0
M1305 8 437 751 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=103710 $D=0
M1306 438 750 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=99080 $D=0
M1307 439 751 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=103710 $D=0
M1308 436 73 438 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=99080 $D=0
M1309 437 73 439 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=103710 $D=0
M1310 438 434 246 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=99080 $D=0
M1311 439 435 247 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=103710 $D=0
M1312 250 440 438 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=99080 $D=0
M1313 251 441 439 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=103710 $D=0
M1314 440 75 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=99080 $D=0
M1315 441 75 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=103710 $D=0
M1316 8 76 442 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=99080 $D=0
M1317 8 76 443 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=103710 $D=0
M1318 444 77 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=99080 $D=0
M1319 445 77 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=103710 $D=0
M1320 446 442 236 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=99080 $D=0
M1321 447 443 237 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=103710 $D=0
M1322 8 446 752 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=99080 $D=0
M1323 8 447 753 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=103710 $D=0
M1324 448 752 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=99080 $D=0
M1325 449 753 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=103710 $D=0
M1326 446 76 448 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=99080 $D=0
M1327 447 76 449 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=103710 $D=0
M1328 448 444 246 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=99080 $D=0
M1329 449 445 247 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=103710 $D=0
M1330 250 450 448 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=99080 $D=0
M1331 251 451 449 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=103710 $D=0
M1332 450 78 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=99080 $D=0
M1333 451 78 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=103710 $D=0
M1334 8 79 452 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=99080 $D=0
M1335 8 79 453 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=103710 $D=0
M1336 454 80 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=99080 $D=0
M1337 455 80 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=103710 $D=0
M1338 456 452 236 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=99080 $D=0
M1339 457 453 237 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=103710 $D=0
M1340 8 456 754 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=99080 $D=0
M1341 8 457 755 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=103710 $D=0
M1342 458 754 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=99080 $D=0
M1343 459 755 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=103710 $D=0
M1344 456 79 458 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=99080 $D=0
M1345 457 79 459 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=103710 $D=0
M1346 458 454 246 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=99080 $D=0
M1347 459 455 247 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=103710 $D=0
M1348 250 460 458 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=99080 $D=0
M1349 251 461 459 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=103710 $D=0
M1350 460 81 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=99080 $D=0
M1351 461 81 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=103710 $D=0
M1352 8 82 462 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=99080 $D=0
M1353 8 82 463 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=103710 $D=0
M1354 464 83 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=99080 $D=0
M1355 465 83 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=103710 $D=0
M1356 466 462 236 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=99080 $D=0
M1357 467 463 237 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=103710 $D=0
M1358 8 466 756 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=99080 $D=0
M1359 8 467 757 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=103710 $D=0
M1360 468 756 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=99080 $D=0
M1361 469 757 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=103710 $D=0
M1362 466 82 468 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=99080 $D=0
M1363 467 82 469 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=103710 $D=0
M1364 468 464 246 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=99080 $D=0
M1365 469 465 247 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=103710 $D=0
M1366 250 470 468 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=99080 $D=0
M1367 251 471 469 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=103710 $D=0
M1368 470 84 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=99080 $D=0
M1369 471 84 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=103710 $D=0
M1370 8 85 472 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=99080 $D=0
M1371 8 85 473 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=103710 $D=0
M1372 474 86 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=99080 $D=0
M1373 475 86 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=103710 $D=0
M1374 476 472 236 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=99080 $D=0
M1375 477 473 237 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=103710 $D=0
M1376 8 476 758 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=99080 $D=0
M1377 8 477 759 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=103710 $D=0
M1378 478 758 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=99080 $D=0
M1379 479 759 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=103710 $D=0
M1380 476 85 478 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=99080 $D=0
M1381 477 85 479 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=103710 $D=0
M1382 478 474 246 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=99080 $D=0
M1383 479 475 247 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=103710 $D=0
M1384 250 480 478 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=99080 $D=0
M1385 251 481 479 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=103710 $D=0
M1386 480 87 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=99080 $D=0
M1387 481 87 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=103710 $D=0
M1388 8 88 482 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=99080 $D=0
M1389 8 88 483 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=103710 $D=0
M1390 484 89 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=99080 $D=0
M1391 485 89 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=103710 $D=0
M1392 486 482 236 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=99080 $D=0
M1393 487 483 237 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=103710 $D=0
M1394 8 486 760 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=99080 $D=0
M1395 8 487 761 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=103710 $D=0
M1396 488 760 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=99080 $D=0
M1397 489 761 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=103710 $D=0
M1398 486 88 488 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=99080 $D=0
M1399 487 88 489 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=103710 $D=0
M1400 488 484 246 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=99080 $D=0
M1401 489 485 247 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=103710 $D=0
M1402 250 490 488 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=99080 $D=0
M1403 251 491 489 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=103710 $D=0
M1404 490 90 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=99080 $D=0
M1405 491 90 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=103710 $D=0
M1406 8 91 492 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=99080 $D=0
M1407 8 91 493 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=103710 $D=0
M1408 494 92 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=99080 $D=0
M1409 495 92 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=103710 $D=0
M1410 496 492 236 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=99080 $D=0
M1411 497 493 237 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=103710 $D=0
M1412 8 496 762 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=99080 $D=0
M1413 8 497 763 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=103710 $D=0
M1414 498 762 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=99080 $D=0
M1415 499 763 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=103710 $D=0
M1416 496 91 498 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=99080 $D=0
M1417 497 91 499 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=103710 $D=0
M1418 498 494 246 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=99080 $D=0
M1419 499 495 247 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=103710 $D=0
M1420 250 500 498 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=99080 $D=0
M1421 251 501 499 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=103710 $D=0
M1422 500 93 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=99080 $D=0
M1423 501 93 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=103710 $D=0
M1424 8 94 502 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=99080 $D=0
M1425 8 94 503 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=103710 $D=0
M1426 504 95 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=99080 $D=0
M1427 505 95 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=103710 $D=0
M1428 506 502 236 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=99080 $D=0
M1429 507 503 237 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=103710 $D=0
M1430 8 506 764 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=99080 $D=0
M1431 8 507 765 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=103710 $D=0
M1432 508 764 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=99080 $D=0
M1433 509 765 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=103710 $D=0
M1434 506 94 508 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=99080 $D=0
M1435 507 94 509 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=103710 $D=0
M1436 508 504 246 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=99080 $D=0
M1437 509 505 247 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=103710 $D=0
M1438 250 510 508 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=99080 $D=0
M1439 251 511 509 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=103710 $D=0
M1440 510 96 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=99080 $D=0
M1441 511 96 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=103710 $D=0
M1442 8 97 512 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=99080 $D=0
M1443 8 97 513 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=103710 $D=0
M1444 514 98 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=99080 $D=0
M1445 515 98 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=103710 $D=0
M1446 516 512 236 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=99080 $D=0
M1447 517 513 237 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=103710 $D=0
M1448 8 516 766 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=99080 $D=0
M1449 8 517 767 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=103710 $D=0
M1450 518 766 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=99080 $D=0
M1451 519 767 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=103710 $D=0
M1452 516 97 518 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=99080 $D=0
M1453 517 97 519 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=103710 $D=0
M1454 518 514 246 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=99080 $D=0
M1455 519 515 247 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=103710 $D=0
M1456 250 520 518 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=99080 $D=0
M1457 251 521 519 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=103710 $D=0
M1458 520 99 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=99080 $D=0
M1459 521 99 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=103710 $D=0
M1460 8 100 522 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=99080 $D=0
M1461 8 100 523 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=103710 $D=0
M1462 524 101 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=99080 $D=0
M1463 525 101 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=103710 $D=0
M1464 526 522 236 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=99080 $D=0
M1465 527 523 237 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=103710 $D=0
M1466 8 526 768 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=99080 $D=0
M1467 8 527 769 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=103710 $D=0
M1468 528 768 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=99080 $D=0
M1469 529 769 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=103710 $D=0
M1470 526 100 528 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=99080 $D=0
M1471 527 100 529 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=103710 $D=0
M1472 528 524 246 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=99080 $D=0
M1473 529 525 247 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=103710 $D=0
M1474 250 530 528 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=99080 $D=0
M1475 251 531 529 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=103710 $D=0
M1476 530 102 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=99080 $D=0
M1477 531 102 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=103710 $D=0
M1478 8 103 532 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=99080 $D=0
M1479 8 103 533 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=103710 $D=0
M1480 534 104 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=99080 $D=0
M1481 535 104 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=103710 $D=0
M1482 536 532 236 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=99080 $D=0
M1483 537 533 237 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=103710 $D=0
M1484 8 536 770 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=99080 $D=0
M1485 8 537 771 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=103710 $D=0
M1486 538 770 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=99080 $D=0
M1487 539 771 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=103710 $D=0
M1488 536 103 538 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=99080 $D=0
M1489 537 103 539 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=103710 $D=0
M1490 538 534 246 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=99080 $D=0
M1491 539 535 247 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=103710 $D=0
M1492 250 540 538 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=99080 $D=0
M1493 251 541 539 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=103710 $D=0
M1494 540 105 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=99080 $D=0
M1495 541 105 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=103710 $D=0
M1496 8 106 542 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=99080 $D=0
M1497 8 106 543 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=103710 $D=0
M1498 544 107 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=99080 $D=0
M1499 545 107 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=103710 $D=0
M1500 546 542 236 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=99080 $D=0
M1501 547 543 237 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=103710 $D=0
M1502 8 546 772 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=99080 $D=0
M1503 8 547 773 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=103710 $D=0
M1504 548 772 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=99080 $D=0
M1505 549 773 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=103710 $D=0
M1506 546 106 548 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=99080 $D=0
M1507 547 106 549 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=103710 $D=0
M1508 548 544 246 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=99080 $D=0
M1509 549 545 247 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=103710 $D=0
M1510 250 550 548 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=99080 $D=0
M1511 251 551 549 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=103710 $D=0
M1512 550 108 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=99080 $D=0
M1513 551 108 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=103710 $D=0
M1514 8 109 552 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=99080 $D=0
M1515 8 109 553 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=103710 $D=0
M1516 554 110 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=99080 $D=0
M1517 555 110 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=103710 $D=0
M1518 5 554 246 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=99080 $D=0
M1519 5 555 247 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=103710 $D=0
M1520 250 552 5 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=99080 $D=0
M1521 251 553 5 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=103710 $D=0
M1522 8 558 556 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=99080 $D=0
M1523 8 559 557 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=103710 $D=0
M1524 558 111 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=99080 $D=0
M1525 559 111 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=103710 $D=0
M1526 774 246 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=99080 $D=0
M1527 775 247 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=103710 $D=0
M1528 560 558 774 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=99080 $D=0
M1529 561 559 775 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=103710 $D=0
M1530 8 560 562 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=99080 $D=0
M1531 8 561 563 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=103710 $D=0
M1532 776 562 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=99080 $D=0
M1533 777 563 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=103710 $D=0
M1534 560 556 776 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=99080 $D=0
M1535 561 557 777 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=103710 $D=0
M1536 8 566 564 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=99080 $D=0
M1537 8 567 565 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=103710 $D=0
M1538 566 111 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=99080 $D=0
M1539 567 111 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=103710 $D=0
M1540 778 250 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=99080 $D=0
M1541 779 251 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=103710 $D=0
M1542 568 566 778 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=99080 $D=0
M1543 569 567 779 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=103710 $D=0
M1544 8 568 112 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=99080 $D=0
M1545 8 569 113 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=103710 $D=0
M1546 780 112 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=99080 $D=0
M1547 781 113 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=103710 $D=0
M1548 568 564 780 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=99080 $D=0
M1549 569 565 781 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=103710 $D=0
M1550 570 115 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=99080 $D=0
M1551 571 115 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=103710 $D=0
M1552 572 115 562 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=99080 $D=0
M1553 573 115 563 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=103710 $D=0
M1554 117 570 572 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=99080 $D=0
M1555 118 571 573 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=103710 $D=0
M1556 574 119 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=99080 $D=0
M1557 575 119 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=103710 $D=0
M1558 576 119 112 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=99080 $D=0
M1559 577 119 113 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=103710 $D=0
M1560 782 574 576 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=99080 $D=0
M1561 783 575 577 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=103710 $D=0
M1562 8 112 782 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=99080 $D=0
M1563 8 113 783 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=103710 $D=0
M1564 578 122 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=99080 $D=0
M1565 579 122 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=103710 $D=0
M1566 580 122 576 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=99080 $D=0
M1567 581 122 577 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=103710 $D=0
M1568 10 578 580 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=99080 $D=0
M1569 11 579 581 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=103710 $D=0
M1570 583 582 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=99080 $D=0
M1571 584 123 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=103710 $D=0
M1572 8 587 585 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=99080 $D=0
M1573 8 588 586 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=103710 $D=0
M1574 589 572 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=99080 $D=0
M1575 590 573 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=103710 $D=0
M1576 587 572 582 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=99080 $D=0
M1577 588 573 123 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=103710 $D=0
M1578 583 589 587 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=99080 $D=0
M1579 584 590 588 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=103710 $D=0
M1580 591 585 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=99080 $D=0
M1581 592 586 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=103710 $D=0
M1582 126 585 580 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=99080 $D=0
M1583 582 586 581 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=103710 $D=0
M1584 572 591 126 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=99080 $D=0
M1585 573 592 582 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=103710 $D=0
M1586 593 126 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=99080 $D=0
M1587 594 582 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=103710 $D=0
M1588 595 585 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=99080 $D=0
M1589 596 586 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=103710 $D=0
M1590 597 585 593 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=99080 $D=0
M1591 598 586 594 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=103710 $D=0
M1592 580 595 597 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=99080 $D=0
M1593 581 596 598 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=103710 $D=0
M1594 794 572 8 8 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=98720 $D=0
M1595 795 573 8 8 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=103350 $D=0
M1596 599 580 794 8 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=98720 $D=0
M1597 600 581 795 8 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=103350 $D=0
M1598 601 597 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=99080 $D=0
M1599 602 598 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=103710 $D=0
M1600 603 572 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=99080 $D=0
M1601 604 573 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=103710 $D=0
M1602 8 580 603 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=99080 $D=0
M1603 8 581 604 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=103710 $D=0
M1604 605 572 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=99080 $D=0
M1605 606 573 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=103710 $D=0
M1606 8 580 605 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=99080 $D=0
M1607 8 581 606 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=103710 $D=0
M1608 796 572 8 8 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=98900 $D=0
M1609 797 573 8 8 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=103530 $D=0
M1610 609 580 796 8 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=98900 $D=0
M1611 610 581 797 8 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=103530 $D=0
M1612 8 605 609 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=99080 $D=0
M1613 8 606 610 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=103710 $D=0
M1614 611 128 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=99080 $D=0
M1615 612 128 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=103710 $D=0
M1616 613 128 599 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=99080 $D=0
M1617 614 128 600 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=103710 $D=0
M1618 603 611 613 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=99080 $D=0
M1619 604 612 614 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=103710 $D=0
M1620 615 128 601 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=99080 $D=0
M1621 616 128 602 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=103710 $D=0
M1622 609 611 615 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=99080 $D=0
M1623 610 612 616 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=103710 $D=0
M1624 617 129 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=99080 $D=0
M1625 618 129 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=103710 $D=0
M1626 619 129 615 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=99080 $D=0
M1627 620 129 616 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=103710 $D=0
M1628 613 617 619 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=99080 $D=0
M1629 614 618 620 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=103710 $D=0
M1630 12 619 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=99080 $D=0
M1631 13 620 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=103710 $D=0
M1632 621 130 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=99080 $D=0
M1633 622 130 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=103710 $D=0
M1634 623 130 131 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=99080 $D=0
M1635 624 130 132 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=103710 $D=0
M1636 133 621 623 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=99080 $D=0
M1637 134 622 624 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=103710 $D=0
M1638 625 130 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=99080 $D=0
M1639 626 130 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=103710 $D=0
M1640 627 130 135 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=99080 $D=0
M1641 628 130 136 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=103710 $D=0
M1642 137 625 627 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=99080 $D=0
M1643 138 626 628 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=103710 $D=0
M1644 629 130 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=99080 $D=0
M1645 630 130 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=103710 $D=0
M1646 631 130 139 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=99080 $D=0
M1647 632 130 140 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=103710 $D=0
M1648 116 629 631 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=99080 $D=0
M1649 121 630 632 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=103710 $D=0
M1650 633 130 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=99080 $D=0
M1651 634 130 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=103710 $D=0
M1652 635 130 141 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=99080 $D=0
M1653 636 130 142 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=103710 $D=0
M1654 114 633 635 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=99080 $D=0
M1655 120 634 636 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=103710 $D=0
M1656 637 130 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=99080 $D=0
M1657 638 130 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=103710 $D=0
M1658 639 130 5 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=99080 $D=0
M1659 640 130 5 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=103710 $D=0
M1660 143 637 639 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=99080 $D=0
M1661 144 638 640 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=103710 $D=0
M1662 8 572 784 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=99080 $D=0
M1663 8 573 785 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=103710 $D=0
M1664 134 784 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=99080 $D=0
M1665 131 785 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=103710 $D=0
M1666 641 145 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=99080 $D=0
M1667 642 145 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=103710 $D=0
M1668 146 145 134 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=99080 $D=0
M1669 147 145 131 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=103710 $D=0
M1670 623 641 146 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=99080 $D=0
M1671 624 642 147 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=103710 $D=0
M1672 643 148 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=99080 $D=0
M1673 644 148 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=103710 $D=0
M1674 149 148 146 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=99080 $D=0
M1675 127 148 147 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=103710 $D=0
M1676 627 643 149 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=99080 $D=0
M1677 628 644 127 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=103710 $D=0
M1678 645 150 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=99080 $D=0
M1679 646 150 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=103710 $D=0
M1680 124 150 149 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=99080 $D=0
M1681 125 150 127 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=103710 $D=0
M1682 631 645 124 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=99080 $D=0
M1683 632 646 125 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=103710 $D=0
M1684 647 151 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=99080 $D=0
M1685 648 151 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=103710 $D=0
M1686 152 151 124 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=99080 $D=0
M1687 153 151 125 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=103710 $D=0
M1688 635 647 152 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=99080 $D=0
M1689 636 648 153 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=103710 $D=0
M1690 649 154 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=99080 $D=0
M1691 650 154 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=103710 $D=0
M1692 222 154 152 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=99080 $D=0
M1693 223 154 153 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=103710 $D=0
M1694 639 649 222 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=99080 $D=0
M1695 640 650 223 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=103710 $D=0
M1696 651 155 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=99080 $D=0
M1697 652 155 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=103710 $D=0
M1698 653 155 112 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=99080 $D=0
M1699 654 155 113 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=103710 $D=0
M1700 10 651 653 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=99080 $D=0
M1701 11 652 654 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=103710 $D=0
M1702 655 562 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=99080 $D=0
M1703 656 563 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=103710 $D=0
M1704 8 653 655 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=99080 $D=0
M1705 8 654 656 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=103710 $D=0
M1706 798 562 8 8 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=98900 $D=0
M1707 799 563 8 8 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=103530 $D=0
M1708 659 653 798 8 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=98900 $D=0
M1709 660 654 799 8 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=103530 $D=0
M1710 8 655 659 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=99080 $D=0
M1711 8 656 660 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=103710 $D=0
M1712 786 156 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=99080 $D=0
M1713 787 661 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=103710 $D=0
M1714 8 659 786 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=99080 $D=0
M1715 8 660 787 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=103710 $D=0
M1716 661 786 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=99080 $D=0
M1717 157 787 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=103710 $D=0
M1718 800 562 8 8 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=98720 $D=0
M1719 801 563 8 8 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=103350 $D=0
M1720 662 664 800 8 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=98720 $D=0
M1721 663 665 801 8 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=103350 $D=0
M1722 664 653 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=99080 $D=0
M1723 665 654 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=103710 $D=0
M1724 666 662 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=99080 $D=0
M1725 667 663 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=103710 $D=0
M1726 8 156 666 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=99080 $D=0
M1727 8 661 667 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=103710 $D=0
M1728 669 158 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=99080 $D=0
M1729 670 668 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=103710 $D=0
M1730 668 666 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=99080 $D=0
M1731 159 667 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=103710 $D=0
M1732 8 669 668 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=99080 $D=0
M1733 8 670 159 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=103710 $D=0
M1734 672 671 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=99080 $D=0
M1735 673 160 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=103710 $D=0
M1736 8 676 674 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=99080 $D=0
M1737 8 677 675 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=103710 $D=0
M1738 678 117 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=99080 $D=0
M1739 679 118 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=103710 $D=0
M1740 676 117 671 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=99080 $D=0
M1741 677 118 160 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=103710 $D=0
M1742 672 678 676 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=99080 $D=0
M1743 673 679 677 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=103710 $D=0
M1744 680 674 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=99080 $D=0
M1745 681 675 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=103710 $D=0
M1746 161 674 5 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=99080 $D=0
M1747 671 675 5 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=103710 $D=0
M1748 117 680 161 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=99080 $D=0
M1749 118 681 671 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=103710 $D=0
M1750 682 161 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=99080 $D=0
M1751 683 671 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=103710 $D=0
M1752 684 674 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=99080 $D=0
M1753 685 675 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=103710 $D=0
M1754 224 674 682 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=99080 $D=0
M1755 225 675 683 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=103710 $D=0
M1756 5 684 224 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=99080 $D=0
M1757 5 685 225 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=103710 $D=0
M1758 686 162 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=99080 $D=0
M1759 687 162 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=103710 $D=0
M1760 688 162 224 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=99080 $D=0
M1761 689 162 225 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=103710 $D=0
M1762 12 686 688 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=99080 $D=0
M1763 13 687 689 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=103710 $D=0
M1764 690 163 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=99080 $D=0
M1765 691 163 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=103710 $D=0
M1766 692 163 688 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=99080 $D=0
M1767 693 163 689 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=103710 $D=0
M1768 5 690 692 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=99080 $D=0
M1769 5 691 693 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=103710 $D=0
M1770 694 111 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=99080 $D=0
M1771 695 111 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=103710 $D=0
M1772 8 694 696 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=99080 $D=0
M1773 8 695 697 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=103710 $D=0
M1774 698 111 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=99080 $D=0
M1775 699 111 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=103710 $D=0
M1776 700 696 692 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=99080 $D=0
M1777 701 697 693 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=103710 $D=0
M1778 8 700 788 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=99080 $D=0
M1779 8 701 789 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=103710 $D=0
M1780 702 788 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=99080 $D=0
M1781 703 789 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=103710 $D=0
M1782 700 694 702 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=99080 $D=0
M1783 701 695 703 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=103710 $D=0
M1784 704 698 702 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=99080 $D=0
M1785 705 699 703 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=103710 $D=0
M1786 8 708 706 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=99080 $D=0
M1787 8 709 707 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=103710 $D=0
M1788 708 111 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=99080 $D=0
M1789 709 111 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=103710 $D=0
M1790 790 704 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=99080 $D=0
M1791 791 705 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=103710 $D=0
M1792 710 708 790 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=99080 $D=0
M1793 711 709 791 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=103710 $D=0
M1794 8 710 117 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=99080 $D=0
M1795 8 711 118 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=103710 $D=0
M1796 792 117 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=99080 $D=0
M1797 793 118 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=103710 $D=0
M1798 710 706 792 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=99080 $D=0
M1799 711 707 793 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=103710 $D=0
.ENDS
***************************************
.SUBCKT ICV_29 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163
** N=817 EP=163 IP=1514 FDC=1800
M0 202 1 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=88570 $D=1
M1 203 1 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=93200 $D=1
M2 204 202 2 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=88570 $D=1
M3 205 203 3 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=93200 $D=1
M4 5 1 204 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=88570 $D=1
M5 5 1 205 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=93200 $D=1
M6 206 202 4 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=88570 $D=1
M7 207 203 4 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=93200 $D=1
M8 2 1 206 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=88570 $D=1
M9 3 1 207 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=93200 $D=1
M10 208 202 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=88570 $D=1
M11 209 203 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=93200 $D=1
M12 2 1 208 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=88570 $D=1
M13 3 1 209 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=93200 $D=1
M14 212 210 208 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=88570 $D=1
M15 213 211 209 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=93200 $D=1
M16 210 6 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=88570 $D=1
M17 211 6 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=93200 $D=1
M18 214 210 206 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=88570 $D=1
M19 215 211 207 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=93200 $D=1
M20 204 6 214 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=88570 $D=1
M21 205 6 215 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=93200 $D=1
M22 216 7 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=88570 $D=1
M23 217 7 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=93200 $D=1
M24 218 216 214 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=88570 $D=1
M25 219 217 215 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=93200 $D=1
M26 212 7 218 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=88570 $D=1
M27 213 7 219 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=93200 $D=1
M28 220 9 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=88570 $D=1
M29 221 9 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=93200 $D=1
M30 222 220 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=88570 $D=1
M31 223 221 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=93200 $D=1
M32 10 9 222 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=88570 $D=1
M33 11 9 223 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=93200 $D=1
M34 224 220 12 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=88570 $D=1
M35 225 221 13 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=93200 $D=1
M36 226 9 224 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=88570 $D=1
M37 227 9 225 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=93200 $D=1
M38 230 220 228 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=88570 $D=1
M39 231 221 229 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=93200 $D=1
M40 218 9 230 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=88570 $D=1
M41 219 9 231 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=93200 $D=1
M42 234 232 230 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=88570 $D=1
M43 235 233 231 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=93200 $D=1
M44 232 14 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=88570 $D=1
M45 233 14 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=93200 $D=1
M46 236 232 224 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=88570 $D=1
M47 237 233 225 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=93200 $D=1
M48 222 14 236 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=88570 $D=1
M49 223 14 237 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=93200 $D=1
M50 238 15 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=88570 $D=1
M51 239 15 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=93200 $D=1
M52 240 238 236 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=88570 $D=1
M53 241 239 237 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=93200 $D=1
M54 234 15 240 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=88570 $D=1
M55 235 15 241 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=93200 $D=1
M56 5 16 242 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=88570 $D=1
M57 5 16 243 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=93200 $D=1
M58 244 17 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=88570 $D=1
M59 245 17 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=93200 $D=1
M60 246 16 240 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=88570 $D=1
M61 247 16 241 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=93200 $D=1
M62 5 246 716 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=88570 $D=1
M63 5 247 717 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=93200 $D=1
M64 248 716 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=88570 $D=1
M65 249 717 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=93200 $D=1
M66 246 242 248 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=88570 $D=1
M67 247 243 249 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=93200 $D=1
M68 248 17 250 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=88570 $D=1
M69 249 17 251 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=93200 $D=1
M70 254 18 248 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=88570 $D=1
M71 255 18 249 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=93200 $D=1
M72 252 18 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=88570 $D=1
M73 253 18 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=93200 $D=1
M74 5 19 256 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=88570 $D=1
M75 5 19 257 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=93200 $D=1
M76 258 20 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=88570 $D=1
M77 259 20 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=93200 $D=1
M78 260 19 240 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=88570 $D=1
M79 261 19 241 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=93200 $D=1
M80 5 260 718 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=88570 $D=1
M81 5 261 719 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=93200 $D=1
M82 262 718 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=88570 $D=1
M83 263 719 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=93200 $D=1
M84 260 256 262 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=88570 $D=1
M85 261 257 263 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=93200 $D=1
M86 262 20 250 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=88570 $D=1
M87 263 20 251 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=93200 $D=1
M88 254 21 262 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=88570 $D=1
M89 255 21 263 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=93200 $D=1
M90 264 21 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=88570 $D=1
M91 265 21 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=93200 $D=1
M92 5 22 266 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=88570 $D=1
M93 5 22 267 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=93200 $D=1
M94 268 23 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=88570 $D=1
M95 269 23 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=93200 $D=1
M96 270 22 240 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=88570 $D=1
M97 271 22 241 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=93200 $D=1
M98 5 270 720 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=88570 $D=1
M99 5 271 721 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=93200 $D=1
M100 272 720 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=88570 $D=1
M101 273 721 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=93200 $D=1
M102 270 266 272 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=88570 $D=1
M103 271 267 273 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=93200 $D=1
M104 272 23 250 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=88570 $D=1
M105 273 23 251 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=93200 $D=1
M106 254 24 272 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=88570 $D=1
M107 255 24 273 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=93200 $D=1
M108 274 24 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=88570 $D=1
M109 275 24 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=93200 $D=1
M110 5 25 276 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=88570 $D=1
M111 5 25 277 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=93200 $D=1
M112 278 26 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=88570 $D=1
M113 279 26 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=93200 $D=1
M114 280 25 240 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=88570 $D=1
M115 281 25 241 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=93200 $D=1
M116 5 280 722 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=88570 $D=1
M117 5 281 723 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=93200 $D=1
M118 282 722 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=88570 $D=1
M119 283 723 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=93200 $D=1
M120 280 276 282 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=88570 $D=1
M121 281 277 283 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=93200 $D=1
M122 282 26 250 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=88570 $D=1
M123 283 26 251 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=93200 $D=1
M124 254 27 282 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=88570 $D=1
M125 255 27 283 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=93200 $D=1
M126 284 27 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=88570 $D=1
M127 285 27 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=93200 $D=1
M128 5 28 286 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=88570 $D=1
M129 5 28 287 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=93200 $D=1
M130 288 29 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=88570 $D=1
M131 289 29 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=93200 $D=1
M132 290 28 240 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=88570 $D=1
M133 291 28 241 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=93200 $D=1
M134 5 290 724 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=88570 $D=1
M135 5 291 725 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=93200 $D=1
M136 292 724 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=88570 $D=1
M137 293 725 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=93200 $D=1
M138 290 286 292 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=88570 $D=1
M139 291 287 293 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=93200 $D=1
M140 292 29 250 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=88570 $D=1
M141 293 29 251 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=93200 $D=1
M142 254 30 292 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=88570 $D=1
M143 255 30 293 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=93200 $D=1
M144 294 30 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=88570 $D=1
M145 295 30 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=93200 $D=1
M146 5 31 296 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=88570 $D=1
M147 5 31 297 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=93200 $D=1
M148 298 32 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=88570 $D=1
M149 299 32 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=93200 $D=1
M150 300 31 240 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=88570 $D=1
M151 301 31 241 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=93200 $D=1
M152 5 300 726 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=88570 $D=1
M153 5 301 727 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=93200 $D=1
M154 302 726 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=88570 $D=1
M155 303 727 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=93200 $D=1
M156 300 296 302 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=88570 $D=1
M157 301 297 303 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=93200 $D=1
M158 302 32 250 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=88570 $D=1
M159 303 32 251 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=93200 $D=1
M160 254 33 302 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=88570 $D=1
M161 255 33 303 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=93200 $D=1
M162 304 33 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=88570 $D=1
M163 305 33 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=93200 $D=1
M164 5 34 306 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=88570 $D=1
M165 5 34 307 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=93200 $D=1
M166 308 35 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=88570 $D=1
M167 309 35 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=93200 $D=1
M168 310 34 240 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=88570 $D=1
M169 311 34 241 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=93200 $D=1
M170 5 310 728 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=88570 $D=1
M171 5 311 729 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=93200 $D=1
M172 312 728 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=88570 $D=1
M173 313 729 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=93200 $D=1
M174 310 306 312 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=88570 $D=1
M175 311 307 313 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=93200 $D=1
M176 312 35 250 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=88570 $D=1
M177 313 35 251 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=93200 $D=1
M178 254 36 312 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=88570 $D=1
M179 255 36 313 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=93200 $D=1
M180 314 36 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=88570 $D=1
M181 315 36 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=93200 $D=1
M182 5 37 316 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=88570 $D=1
M183 5 37 317 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=93200 $D=1
M184 318 38 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=88570 $D=1
M185 319 38 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=93200 $D=1
M186 320 37 240 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=88570 $D=1
M187 321 37 241 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=93200 $D=1
M188 5 320 730 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=88570 $D=1
M189 5 321 731 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=93200 $D=1
M190 322 730 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=88570 $D=1
M191 323 731 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=93200 $D=1
M192 320 316 322 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=88570 $D=1
M193 321 317 323 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=93200 $D=1
M194 322 38 250 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=88570 $D=1
M195 323 38 251 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=93200 $D=1
M196 254 39 322 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=88570 $D=1
M197 255 39 323 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=93200 $D=1
M198 324 39 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=88570 $D=1
M199 325 39 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=93200 $D=1
M200 5 40 326 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=88570 $D=1
M201 5 40 327 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=93200 $D=1
M202 328 41 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=88570 $D=1
M203 329 41 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=93200 $D=1
M204 330 40 240 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=88570 $D=1
M205 331 40 241 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=93200 $D=1
M206 5 330 732 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=88570 $D=1
M207 5 331 733 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=93200 $D=1
M208 332 732 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=88570 $D=1
M209 333 733 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=93200 $D=1
M210 330 326 332 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=88570 $D=1
M211 331 327 333 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=93200 $D=1
M212 332 41 250 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=88570 $D=1
M213 333 41 251 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=93200 $D=1
M214 254 42 332 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=88570 $D=1
M215 255 42 333 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=93200 $D=1
M216 334 42 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=88570 $D=1
M217 335 42 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=93200 $D=1
M218 5 43 336 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=88570 $D=1
M219 5 43 337 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=93200 $D=1
M220 338 44 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=88570 $D=1
M221 339 44 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=93200 $D=1
M222 340 43 240 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=88570 $D=1
M223 341 43 241 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=93200 $D=1
M224 5 340 734 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=88570 $D=1
M225 5 341 735 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=93200 $D=1
M226 342 734 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=88570 $D=1
M227 343 735 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=93200 $D=1
M228 340 336 342 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=88570 $D=1
M229 341 337 343 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=93200 $D=1
M230 342 44 250 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=88570 $D=1
M231 343 44 251 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=93200 $D=1
M232 254 45 342 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=88570 $D=1
M233 255 45 343 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=93200 $D=1
M234 344 45 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=88570 $D=1
M235 345 45 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=93200 $D=1
M236 5 46 346 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=88570 $D=1
M237 5 46 347 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=93200 $D=1
M238 348 47 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=88570 $D=1
M239 349 47 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=93200 $D=1
M240 350 46 240 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=88570 $D=1
M241 351 46 241 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=93200 $D=1
M242 5 350 736 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=88570 $D=1
M243 5 351 737 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=93200 $D=1
M244 352 736 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=88570 $D=1
M245 353 737 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=93200 $D=1
M246 350 346 352 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=88570 $D=1
M247 351 347 353 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=93200 $D=1
M248 352 47 250 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=88570 $D=1
M249 353 47 251 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=93200 $D=1
M250 254 48 352 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=88570 $D=1
M251 255 48 353 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=93200 $D=1
M252 354 48 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=88570 $D=1
M253 355 48 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=93200 $D=1
M254 5 49 356 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=88570 $D=1
M255 5 49 357 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=93200 $D=1
M256 358 50 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=88570 $D=1
M257 359 50 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=93200 $D=1
M258 360 49 240 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=88570 $D=1
M259 361 49 241 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=93200 $D=1
M260 5 360 738 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=88570 $D=1
M261 5 361 739 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=93200 $D=1
M262 362 738 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=88570 $D=1
M263 363 739 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=93200 $D=1
M264 360 356 362 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=88570 $D=1
M265 361 357 363 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=93200 $D=1
M266 362 50 250 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=88570 $D=1
M267 363 50 251 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=93200 $D=1
M268 254 51 362 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=88570 $D=1
M269 255 51 363 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=93200 $D=1
M270 364 51 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=88570 $D=1
M271 365 51 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=93200 $D=1
M272 5 52 366 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=88570 $D=1
M273 5 52 367 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=93200 $D=1
M274 368 53 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=88570 $D=1
M275 369 53 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=93200 $D=1
M276 370 52 240 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=88570 $D=1
M277 371 52 241 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=93200 $D=1
M278 5 370 740 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=88570 $D=1
M279 5 371 741 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=93200 $D=1
M280 372 740 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=88570 $D=1
M281 373 741 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=93200 $D=1
M282 370 366 372 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=88570 $D=1
M283 371 367 373 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=93200 $D=1
M284 372 53 250 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=88570 $D=1
M285 373 53 251 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=93200 $D=1
M286 254 54 372 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=88570 $D=1
M287 255 54 373 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=93200 $D=1
M288 374 54 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=88570 $D=1
M289 375 54 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=93200 $D=1
M290 5 55 376 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=88570 $D=1
M291 5 55 377 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=93200 $D=1
M292 378 56 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=88570 $D=1
M293 379 56 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=93200 $D=1
M294 380 55 240 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=88570 $D=1
M295 381 55 241 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=93200 $D=1
M296 5 380 742 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=88570 $D=1
M297 5 381 743 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=93200 $D=1
M298 382 742 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=88570 $D=1
M299 383 743 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=93200 $D=1
M300 380 376 382 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=88570 $D=1
M301 381 377 383 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=93200 $D=1
M302 382 56 250 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=88570 $D=1
M303 383 56 251 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=93200 $D=1
M304 254 57 382 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=88570 $D=1
M305 255 57 383 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=93200 $D=1
M306 384 57 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=88570 $D=1
M307 385 57 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=93200 $D=1
M308 5 58 386 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=88570 $D=1
M309 5 58 387 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=93200 $D=1
M310 388 59 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=88570 $D=1
M311 389 59 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=93200 $D=1
M312 390 58 240 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=88570 $D=1
M313 391 58 241 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=93200 $D=1
M314 5 390 744 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=88570 $D=1
M315 5 391 745 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=93200 $D=1
M316 392 744 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=88570 $D=1
M317 393 745 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=93200 $D=1
M318 390 386 392 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=88570 $D=1
M319 391 387 393 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=93200 $D=1
M320 392 59 250 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=88570 $D=1
M321 393 59 251 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=93200 $D=1
M322 254 60 392 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=88570 $D=1
M323 255 60 393 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=93200 $D=1
M324 394 60 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=88570 $D=1
M325 395 60 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=93200 $D=1
M326 5 61 396 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=88570 $D=1
M327 5 61 397 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=93200 $D=1
M328 398 62 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=88570 $D=1
M329 399 62 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=93200 $D=1
M330 400 61 240 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=88570 $D=1
M331 401 61 241 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=93200 $D=1
M332 5 400 746 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=88570 $D=1
M333 5 401 747 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=93200 $D=1
M334 402 746 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=88570 $D=1
M335 403 747 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=93200 $D=1
M336 400 396 402 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=88570 $D=1
M337 401 397 403 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=93200 $D=1
M338 402 62 250 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=88570 $D=1
M339 403 62 251 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=93200 $D=1
M340 254 63 402 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=88570 $D=1
M341 255 63 403 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=93200 $D=1
M342 404 63 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=88570 $D=1
M343 405 63 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=93200 $D=1
M344 5 64 406 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=88570 $D=1
M345 5 64 407 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=93200 $D=1
M346 408 65 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=88570 $D=1
M347 409 65 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=93200 $D=1
M348 410 64 240 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=88570 $D=1
M349 411 64 241 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=93200 $D=1
M350 5 410 748 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=88570 $D=1
M351 5 411 749 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=93200 $D=1
M352 412 748 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=88570 $D=1
M353 413 749 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=93200 $D=1
M354 410 406 412 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=88570 $D=1
M355 411 407 413 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=93200 $D=1
M356 412 65 250 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=88570 $D=1
M357 413 65 251 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=93200 $D=1
M358 254 66 412 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=88570 $D=1
M359 255 66 413 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=93200 $D=1
M360 414 66 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=88570 $D=1
M361 415 66 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=93200 $D=1
M362 5 67 416 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=88570 $D=1
M363 5 67 417 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=93200 $D=1
M364 418 68 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=88570 $D=1
M365 419 68 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=93200 $D=1
M366 420 67 240 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=88570 $D=1
M367 421 67 241 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=93200 $D=1
M368 5 420 750 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=88570 $D=1
M369 5 421 751 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=93200 $D=1
M370 422 750 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=88570 $D=1
M371 423 751 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=93200 $D=1
M372 420 416 422 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=88570 $D=1
M373 421 417 423 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=93200 $D=1
M374 422 68 250 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=88570 $D=1
M375 423 68 251 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=93200 $D=1
M376 254 69 422 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=88570 $D=1
M377 255 69 423 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=93200 $D=1
M378 424 69 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=88570 $D=1
M379 425 69 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=93200 $D=1
M380 5 70 426 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=88570 $D=1
M381 5 70 427 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=93200 $D=1
M382 428 71 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=88570 $D=1
M383 429 71 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=93200 $D=1
M384 430 70 240 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=88570 $D=1
M385 431 70 241 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=93200 $D=1
M386 5 430 752 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=88570 $D=1
M387 5 431 753 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=93200 $D=1
M388 432 752 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=88570 $D=1
M389 433 753 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=93200 $D=1
M390 430 426 432 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=88570 $D=1
M391 431 427 433 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=93200 $D=1
M392 432 71 250 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=88570 $D=1
M393 433 71 251 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=93200 $D=1
M394 254 72 432 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=88570 $D=1
M395 255 72 433 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=93200 $D=1
M396 434 72 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=88570 $D=1
M397 435 72 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=93200 $D=1
M398 5 73 436 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=88570 $D=1
M399 5 73 437 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=93200 $D=1
M400 438 74 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=88570 $D=1
M401 439 74 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=93200 $D=1
M402 440 73 240 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=88570 $D=1
M403 441 73 241 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=93200 $D=1
M404 5 440 754 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=88570 $D=1
M405 5 441 755 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=93200 $D=1
M406 442 754 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=88570 $D=1
M407 443 755 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=93200 $D=1
M408 440 436 442 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=88570 $D=1
M409 441 437 443 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=93200 $D=1
M410 442 74 250 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=88570 $D=1
M411 443 74 251 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=93200 $D=1
M412 254 75 442 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=88570 $D=1
M413 255 75 443 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=93200 $D=1
M414 444 75 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=88570 $D=1
M415 445 75 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=93200 $D=1
M416 5 76 446 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=88570 $D=1
M417 5 76 447 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=93200 $D=1
M418 448 77 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=88570 $D=1
M419 449 77 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=93200 $D=1
M420 450 76 240 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=88570 $D=1
M421 451 76 241 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=93200 $D=1
M422 5 450 756 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=88570 $D=1
M423 5 451 757 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=93200 $D=1
M424 452 756 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=88570 $D=1
M425 453 757 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=93200 $D=1
M426 450 446 452 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=88570 $D=1
M427 451 447 453 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=93200 $D=1
M428 452 77 250 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=88570 $D=1
M429 453 77 251 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=93200 $D=1
M430 254 78 452 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=88570 $D=1
M431 255 78 453 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=93200 $D=1
M432 454 78 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=88570 $D=1
M433 455 78 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=93200 $D=1
M434 5 79 456 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=88570 $D=1
M435 5 79 457 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=93200 $D=1
M436 458 80 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=88570 $D=1
M437 459 80 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=93200 $D=1
M438 460 79 240 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=88570 $D=1
M439 461 79 241 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=93200 $D=1
M440 5 460 758 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=88570 $D=1
M441 5 461 759 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=93200 $D=1
M442 462 758 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=88570 $D=1
M443 463 759 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=93200 $D=1
M444 460 456 462 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=88570 $D=1
M445 461 457 463 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=93200 $D=1
M446 462 80 250 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=88570 $D=1
M447 463 80 251 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=93200 $D=1
M448 254 81 462 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=88570 $D=1
M449 255 81 463 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=93200 $D=1
M450 464 81 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=88570 $D=1
M451 465 81 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=93200 $D=1
M452 5 82 466 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=88570 $D=1
M453 5 82 467 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=93200 $D=1
M454 468 83 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=88570 $D=1
M455 469 83 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=93200 $D=1
M456 470 82 240 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=88570 $D=1
M457 471 82 241 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=93200 $D=1
M458 5 470 760 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=88570 $D=1
M459 5 471 761 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=93200 $D=1
M460 472 760 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=88570 $D=1
M461 473 761 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=93200 $D=1
M462 470 466 472 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=88570 $D=1
M463 471 467 473 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=93200 $D=1
M464 472 83 250 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=88570 $D=1
M465 473 83 251 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=93200 $D=1
M466 254 84 472 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=88570 $D=1
M467 255 84 473 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=93200 $D=1
M468 474 84 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=88570 $D=1
M469 475 84 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=93200 $D=1
M470 5 85 476 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=88570 $D=1
M471 5 85 477 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=93200 $D=1
M472 478 86 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=88570 $D=1
M473 479 86 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=93200 $D=1
M474 480 85 240 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=88570 $D=1
M475 481 85 241 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=93200 $D=1
M476 5 480 762 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=88570 $D=1
M477 5 481 763 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=93200 $D=1
M478 482 762 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=88570 $D=1
M479 483 763 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=93200 $D=1
M480 480 476 482 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=88570 $D=1
M481 481 477 483 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=93200 $D=1
M482 482 86 250 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=88570 $D=1
M483 483 86 251 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=93200 $D=1
M484 254 87 482 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=88570 $D=1
M485 255 87 483 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=93200 $D=1
M486 484 87 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=88570 $D=1
M487 485 87 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=93200 $D=1
M488 5 88 486 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=88570 $D=1
M489 5 88 487 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=93200 $D=1
M490 488 89 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=88570 $D=1
M491 489 89 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=93200 $D=1
M492 490 88 240 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=88570 $D=1
M493 491 88 241 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=93200 $D=1
M494 5 490 764 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=88570 $D=1
M495 5 491 765 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=93200 $D=1
M496 492 764 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=88570 $D=1
M497 493 765 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=93200 $D=1
M498 490 486 492 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=88570 $D=1
M499 491 487 493 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=93200 $D=1
M500 492 89 250 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=88570 $D=1
M501 493 89 251 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=93200 $D=1
M502 254 90 492 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=88570 $D=1
M503 255 90 493 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=93200 $D=1
M504 494 90 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=88570 $D=1
M505 495 90 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=93200 $D=1
M506 5 91 496 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=88570 $D=1
M507 5 91 497 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=93200 $D=1
M508 498 92 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=88570 $D=1
M509 499 92 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=93200 $D=1
M510 500 91 240 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=88570 $D=1
M511 501 91 241 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=93200 $D=1
M512 5 500 766 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=88570 $D=1
M513 5 501 767 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=93200 $D=1
M514 502 766 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=88570 $D=1
M515 503 767 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=93200 $D=1
M516 500 496 502 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=88570 $D=1
M517 501 497 503 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=93200 $D=1
M518 502 92 250 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=88570 $D=1
M519 503 92 251 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=93200 $D=1
M520 254 93 502 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=88570 $D=1
M521 255 93 503 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=93200 $D=1
M522 504 93 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=88570 $D=1
M523 505 93 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=93200 $D=1
M524 5 94 506 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=88570 $D=1
M525 5 94 507 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=93200 $D=1
M526 508 95 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=88570 $D=1
M527 509 95 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=93200 $D=1
M528 510 94 240 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=88570 $D=1
M529 511 94 241 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=93200 $D=1
M530 5 510 768 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=88570 $D=1
M531 5 511 769 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=93200 $D=1
M532 512 768 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=88570 $D=1
M533 513 769 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=93200 $D=1
M534 510 506 512 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=88570 $D=1
M535 511 507 513 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=93200 $D=1
M536 512 95 250 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=88570 $D=1
M537 513 95 251 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=93200 $D=1
M538 254 96 512 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=88570 $D=1
M539 255 96 513 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=93200 $D=1
M540 514 96 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=88570 $D=1
M541 515 96 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=93200 $D=1
M542 5 97 516 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=88570 $D=1
M543 5 97 517 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=93200 $D=1
M544 518 98 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=88570 $D=1
M545 519 98 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=93200 $D=1
M546 520 97 240 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=88570 $D=1
M547 521 97 241 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=93200 $D=1
M548 5 520 770 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=88570 $D=1
M549 5 521 771 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=93200 $D=1
M550 522 770 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=88570 $D=1
M551 523 771 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=93200 $D=1
M552 520 516 522 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=88570 $D=1
M553 521 517 523 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=93200 $D=1
M554 522 98 250 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=88570 $D=1
M555 523 98 251 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=93200 $D=1
M556 254 99 522 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=88570 $D=1
M557 255 99 523 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=93200 $D=1
M558 524 99 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=88570 $D=1
M559 525 99 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=93200 $D=1
M560 5 100 526 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=88570 $D=1
M561 5 100 527 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=93200 $D=1
M562 528 101 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=88570 $D=1
M563 529 101 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=93200 $D=1
M564 530 100 240 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=88570 $D=1
M565 531 100 241 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=93200 $D=1
M566 5 530 772 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=88570 $D=1
M567 5 531 773 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=93200 $D=1
M568 532 772 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=88570 $D=1
M569 533 773 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=93200 $D=1
M570 530 526 532 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=88570 $D=1
M571 531 527 533 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=93200 $D=1
M572 532 101 250 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=88570 $D=1
M573 533 101 251 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=93200 $D=1
M574 254 102 532 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=88570 $D=1
M575 255 102 533 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=93200 $D=1
M576 534 102 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=88570 $D=1
M577 535 102 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=93200 $D=1
M578 5 103 536 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=88570 $D=1
M579 5 103 537 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=93200 $D=1
M580 538 104 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=88570 $D=1
M581 539 104 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=93200 $D=1
M582 540 103 240 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=88570 $D=1
M583 541 103 241 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=93200 $D=1
M584 5 540 774 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=88570 $D=1
M585 5 541 775 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=93200 $D=1
M586 542 774 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=88570 $D=1
M587 543 775 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=93200 $D=1
M588 540 536 542 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=88570 $D=1
M589 541 537 543 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=93200 $D=1
M590 542 104 250 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=88570 $D=1
M591 543 104 251 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=93200 $D=1
M592 254 105 542 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=88570 $D=1
M593 255 105 543 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=93200 $D=1
M594 544 105 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=88570 $D=1
M595 545 105 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=93200 $D=1
M596 5 106 546 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=88570 $D=1
M597 5 106 547 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=93200 $D=1
M598 548 107 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=88570 $D=1
M599 549 107 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=93200 $D=1
M600 550 106 240 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=88570 $D=1
M601 551 106 241 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=93200 $D=1
M602 5 550 776 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=88570 $D=1
M603 5 551 777 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=93200 $D=1
M604 552 776 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=88570 $D=1
M605 553 777 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=93200 $D=1
M606 550 546 552 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=88570 $D=1
M607 551 547 553 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=93200 $D=1
M608 552 107 250 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=88570 $D=1
M609 553 107 251 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=93200 $D=1
M610 254 108 552 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=88570 $D=1
M611 255 108 553 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=93200 $D=1
M612 554 108 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=88570 $D=1
M613 555 108 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=93200 $D=1
M614 5 109 556 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=88570 $D=1
M615 5 109 557 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=93200 $D=1
M616 558 110 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=88570 $D=1
M617 559 110 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=93200 $D=1
M618 5 110 250 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=88570 $D=1
M619 5 110 251 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=93200 $D=1
M620 254 109 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=88570 $D=1
M621 255 109 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=93200 $D=1
M622 5 562 560 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=88570 $D=1
M623 5 563 561 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=93200 $D=1
M624 562 111 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=88570 $D=1
M625 563 111 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=93200 $D=1
M626 778 250 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=88570 $D=1
M627 779 251 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=93200 $D=1
M628 564 560 778 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=88570 $D=1
M629 565 561 779 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=93200 $D=1
M630 5 564 566 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=88570 $D=1
M631 5 565 567 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=93200 $D=1
M632 780 566 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=88570 $D=1
M633 781 567 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=93200 $D=1
M634 564 562 780 5 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=88570 $D=1
M635 565 563 781 5 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=93200 $D=1
M636 5 570 568 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=88570 $D=1
M637 5 571 569 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=93200 $D=1
M638 570 111 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=88570 $D=1
M639 571 111 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=93200 $D=1
M640 782 254 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=88570 $D=1
M641 783 255 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=93200 $D=1
M642 572 568 782 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=88570 $D=1
M643 573 569 783 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=93200 $D=1
M644 5 572 112 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=88570 $D=1
M645 5 573 113 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=93200 $D=1
M646 784 112 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=88570 $D=1
M647 785 113 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=93200 $D=1
M648 572 570 784 5 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=88570 $D=1
M649 573 571 785 5 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=93200 $D=1
M650 574 118 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=88570 $D=1
M651 575 118 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=93200 $D=1
M652 576 574 566 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=88570 $D=1
M653 577 575 567 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=93200 $D=1
M654 119 118 576 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=88570 $D=1
M655 120 118 577 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=93200 $D=1
M656 578 121 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=88570 $D=1
M657 579 121 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=93200 $D=1
M658 580 578 112 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=88570 $D=1
M659 581 579 113 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=93200 $D=1
M660 786 121 580 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=88570 $D=1
M661 787 121 581 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=93200 $D=1
M662 5 112 786 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=88570 $D=1
M663 5 113 787 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=93200 $D=1
M664 582 123 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=88570 $D=1
M665 583 123 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=93200 $D=1
M666 584 582 580 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=88570 $D=1
M667 585 583 581 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=93200 $D=1
M668 10 123 584 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=88570 $D=1
M669 11 123 585 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=93200 $D=1
M670 587 586 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=88570 $D=1
M671 588 124 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=93200 $D=1
M672 5 591 589 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=88570 $D=1
M673 5 592 590 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=93200 $D=1
M674 593 576 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=88570 $D=1
M675 594 577 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=93200 $D=1
M676 591 593 586 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=88570 $D=1
M677 592 594 124 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=93200 $D=1
M678 587 576 591 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=88570 $D=1
M679 588 577 592 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=93200 $D=1
M680 595 589 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=88570 $D=1
M681 596 590 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=93200 $D=1
M682 127 595 584 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=88570 $D=1
M683 586 596 585 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=93200 $D=1
M684 576 589 127 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=88570 $D=1
M685 577 590 586 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=93200 $D=1
M686 597 127 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=88570 $D=1
M687 598 586 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=93200 $D=1
M688 599 589 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=88570 $D=1
M689 600 590 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=93200 $D=1
M690 601 599 597 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=88570 $D=1
M691 602 600 598 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=93200 $D=1
M692 584 589 601 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=88570 $D=1
M693 585 590 602 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=93200 $D=1
M694 603 576 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=88570 $D=1
M695 604 577 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=93200 $D=1
M696 5 584 603 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=88570 $D=1
M697 5 585 604 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=93200 $D=1
M698 605 601 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=88570 $D=1
M699 606 602 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=93200 $D=1
M700 806 576 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=88570 $D=1
M701 807 577 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=93200 $D=1
M702 607 584 806 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=88570 $D=1
M703 608 585 807 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=93200 $D=1
M704 808 576 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=88570 $D=1
M705 809 577 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=93200 $D=1
M706 609 584 808 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=88570 $D=1
M707 610 585 809 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=93200 $D=1
M708 613 576 611 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=88570 $D=1
M709 614 577 612 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=93200 $D=1
M710 611 584 613 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=88570 $D=1
M711 612 585 614 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=93200 $D=1
M712 5 609 611 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=88570 $D=1
M713 5 610 612 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=93200 $D=1
M714 615 128 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=88570 $D=1
M715 616 128 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=93200 $D=1
M716 617 615 603 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=88570 $D=1
M717 618 616 604 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=93200 $D=1
M718 607 128 617 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=88570 $D=1
M719 608 128 618 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=93200 $D=1
M720 619 615 605 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=88570 $D=1
M721 620 616 606 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=93200 $D=1
M722 613 128 619 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=88570 $D=1
M723 614 128 620 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=93200 $D=1
M724 621 129 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=88570 $D=1
M725 622 129 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=93200 $D=1
M726 623 621 619 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=88570 $D=1
M727 624 622 620 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=93200 $D=1
M728 617 129 623 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=88570 $D=1
M729 618 129 624 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=93200 $D=1
M730 12 623 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=88570 $D=1
M731 13 624 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=93200 $D=1
M732 625 130 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=88570 $D=1
M733 626 130 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=93200 $D=1
M734 627 625 131 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=88570 $D=1
M735 628 626 132 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=93200 $D=1
M736 133 130 627 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=88570 $D=1
M737 134 130 628 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=93200 $D=1
M738 629 130 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=88570 $D=1
M739 630 130 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=93200 $D=1
M740 631 629 135 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=88570 $D=1
M741 632 630 136 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=93200 $D=1
M742 137 130 631 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=88570 $D=1
M743 138 130 632 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=93200 $D=1
M744 633 130 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=88570 $D=1
M745 634 130 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=93200 $D=1
M746 635 633 139 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=88570 $D=1
M747 636 634 140 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=93200 $D=1
M748 114 130 635 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=88570 $D=1
M749 116 130 636 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=93200 $D=1
M750 637 130 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=88570 $D=1
M751 638 130 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=93200 $D=1
M752 639 637 141 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=88570 $D=1
M753 640 638 142 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=93200 $D=1
M754 115 130 639 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=88570 $D=1
M755 117 130 640 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=93200 $D=1
M756 641 130 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=88570 $D=1
M757 642 130 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=93200 $D=1
M758 643 641 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=88570 $D=1
M759 644 642 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=93200 $D=1
M760 143 130 643 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=88570 $D=1
M761 144 130 644 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=93200 $D=1
M762 5 576 788 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=88570 $D=1
M763 5 577 789 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=93200 $D=1
M764 134 788 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=88570 $D=1
M765 131 789 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=93200 $D=1
M766 645 145 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=88570 $D=1
M767 646 145 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=93200 $D=1
M768 146 645 134 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=88570 $D=1
M769 147 646 131 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=93200 $D=1
M770 627 145 146 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=88570 $D=1
M771 628 145 147 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=93200 $D=1
M772 647 148 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=88570 $D=1
M773 648 148 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=93200 $D=1
M774 122 647 146 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=88570 $D=1
M775 149 648 147 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=93200 $D=1
M776 631 148 122 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=88570 $D=1
M777 632 148 149 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=93200 $D=1
M778 649 150 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=88570 $D=1
M779 650 150 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=93200 $D=1
M780 125 649 122 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=88570 $D=1
M781 126 650 149 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=93200 $D=1
M782 635 150 125 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=88570 $D=1
M783 636 150 126 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=93200 $D=1
M784 651 151 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=88570 $D=1
M785 652 151 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=93200 $D=1
M786 152 651 125 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=88570 $D=1
M787 153 652 126 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=93200 $D=1
M788 639 151 152 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=88570 $D=1
M789 640 151 153 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=93200 $D=1
M790 653 154 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=88570 $D=1
M791 654 154 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=93200 $D=1
M792 226 653 152 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=88570 $D=1
M793 227 654 153 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=93200 $D=1
M794 643 154 226 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=88570 $D=1
M795 644 154 227 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=93200 $D=1
M796 655 155 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=88570 $D=1
M797 656 155 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=93200 $D=1
M798 657 655 112 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=88570 $D=1
M799 658 656 113 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=93200 $D=1
M800 10 155 657 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=88570 $D=1
M801 11 155 658 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=93200 $D=1
M802 810 566 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=88570 $D=1
M803 811 567 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=93200 $D=1
M804 659 657 810 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=88570 $D=1
M805 660 658 811 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=93200 $D=1
M806 663 566 661 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=88570 $D=1
M807 664 567 662 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=93200 $D=1
M808 661 657 663 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=88570 $D=1
M809 662 658 664 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=93200 $D=1
M810 5 659 661 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=88570 $D=1
M811 5 660 662 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=93200 $D=1
M812 812 156 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=88570 $D=1
M813 813 665 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=93200 $D=1
M814 790 663 812 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=88570 $D=1
M815 791 664 813 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=93200 $D=1
M816 665 790 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=88570 $D=1
M817 157 791 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=93200 $D=1
M818 666 566 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=88570 $D=1
M819 667 567 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=93200 $D=1
M820 5 668 666 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=88570 $D=1
M821 5 669 667 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=93200 $D=1
M822 668 657 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=88570 $D=1
M823 669 658 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=93200 $D=1
M824 814 666 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=88570 $D=1
M825 815 667 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=93200 $D=1
M826 670 156 814 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=88570 $D=1
M827 671 665 815 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=93200 $D=1
M828 673 158 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=88570 $D=1
M829 674 672 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=93200 $D=1
M830 816 670 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=88570 $D=1
M831 817 671 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=93200 $D=1
M832 672 673 816 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=88570 $D=1
M833 159 674 817 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=93200 $D=1
M834 676 675 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=88570 $D=1
M835 677 160 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=93200 $D=1
M836 5 680 678 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=88570 $D=1
M837 5 681 679 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=93200 $D=1
M838 682 119 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=88570 $D=1
M839 683 120 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=93200 $D=1
M840 680 682 675 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=88570 $D=1
M841 681 683 160 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=93200 $D=1
M842 676 119 680 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=88570 $D=1
M843 677 120 681 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=93200 $D=1
M844 684 678 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=88570 $D=1
M845 685 679 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=93200 $D=1
M846 161 684 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=88570 $D=1
M847 675 685 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=93200 $D=1
M848 119 678 161 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=88570 $D=1
M849 120 679 675 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=93200 $D=1
M850 686 161 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=88570 $D=1
M851 687 675 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=93200 $D=1
M852 688 678 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=88570 $D=1
M853 689 679 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=93200 $D=1
M854 228 688 686 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=88570 $D=1
M855 229 689 687 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=93200 $D=1
M856 5 678 228 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=88570 $D=1
M857 5 679 229 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=93200 $D=1
M858 690 162 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=88570 $D=1
M859 691 162 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=93200 $D=1
M860 692 690 228 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=88570 $D=1
M861 693 691 229 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=93200 $D=1
M862 12 162 692 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=88570 $D=1
M863 13 162 693 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=93200 $D=1
M864 694 163 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=88570 $D=1
M865 695 163 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=93200 $D=1
M866 696 694 692 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=88570 $D=1
M867 697 695 693 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=93200 $D=1
M868 5 163 696 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=88570 $D=1
M869 5 163 697 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=93200 $D=1
M870 698 111 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=88570 $D=1
M871 699 111 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=93200 $D=1
M872 5 698 700 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=88570 $D=1
M873 5 699 701 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=93200 $D=1
M874 702 111 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=88570 $D=1
M875 703 111 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=93200 $D=1
M876 704 698 696 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=88570 $D=1
M877 705 699 697 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=93200 $D=1
M878 5 704 792 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=88570 $D=1
M879 5 705 793 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=93200 $D=1
M880 706 792 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=88570 $D=1
M881 707 793 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=93200 $D=1
M882 704 700 706 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=88570 $D=1
M883 705 701 707 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=93200 $D=1
M884 708 111 706 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=88570 $D=1
M885 709 111 707 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=93200 $D=1
M886 5 712 710 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=88570 $D=1
M887 5 713 711 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=93200 $D=1
M888 712 111 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=88570 $D=1
M889 713 111 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=93200 $D=1
M890 794 708 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=88570 $D=1
M891 795 709 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=93200 $D=1
M892 714 710 794 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=88570 $D=1
M893 715 711 795 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=93200 $D=1
M894 5 714 119 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=88570 $D=1
M895 5 715 120 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=93200 $D=1
M896 796 119 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=88570 $D=1
M897 797 120 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=93200 $D=1
M898 714 712 796 5 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=88570 $D=1
M899 715 713 797 5 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=93200 $D=1
M900 202 1 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=89820 $D=0
M901 203 1 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=94450 $D=0
M902 204 1 2 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=89820 $D=0
M903 205 1 3 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=94450 $D=0
M904 5 202 204 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=89820 $D=0
M905 5 203 205 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=94450 $D=0
M906 206 1 4 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=89820 $D=0
M907 207 1 4 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=94450 $D=0
M908 2 202 206 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=89820 $D=0
M909 3 203 207 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=94450 $D=0
M910 208 1 5 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=89820 $D=0
M911 209 1 5 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=94450 $D=0
M912 2 202 208 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=89820 $D=0
M913 3 203 209 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=94450 $D=0
M914 212 6 208 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=89820 $D=0
M915 213 6 209 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=94450 $D=0
M916 210 6 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=89820 $D=0
M917 211 6 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=94450 $D=0
M918 214 6 206 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=89820 $D=0
M919 215 6 207 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=94450 $D=0
M920 204 210 214 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=89820 $D=0
M921 205 211 215 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=94450 $D=0
M922 216 7 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=89820 $D=0
M923 217 7 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=94450 $D=0
M924 218 7 214 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=89820 $D=0
M925 219 7 215 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=94450 $D=0
M926 212 216 218 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=89820 $D=0
M927 213 217 219 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=94450 $D=0
M928 220 9 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=89820 $D=0
M929 221 9 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=94450 $D=0
M930 222 9 5 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=89820 $D=0
M931 223 9 5 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=94450 $D=0
M932 10 220 222 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=89820 $D=0
M933 11 221 223 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=94450 $D=0
M934 224 9 12 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=89820 $D=0
M935 225 9 13 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=94450 $D=0
M936 226 220 224 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=89820 $D=0
M937 227 221 225 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=94450 $D=0
M938 230 9 228 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=89820 $D=0
M939 231 9 229 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=94450 $D=0
M940 218 220 230 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=89820 $D=0
M941 219 221 231 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=94450 $D=0
M942 234 14 230 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=89820 $D=0
M943 235 14 231 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=94450 $D=0
M944 232 14 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=89820 $D=0
M945 233 14 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=94450 $D=0
M946 236 14 224 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=89820 $D=0
M947 237 14 225 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=94450 $D=0
M948 222 232 236 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=89820 $D=0
M949 223 233 237 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=94450 $D=0
M950 238 15 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=89820 $D=0
M951 239 15 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=94450 $D=0
M952 240 15 236 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=89820 $D=0
M953 241 15 237 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=94450 $D=0
M954 234 238 240 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=89820 $D=0
M955 235 239 241 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=94450 $D=0
M956 8 16 242 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=89820 $D=0
M957 8 16 243 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=94450 $D=0
M958 244 17 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=89820 $D=0
M959 245 17 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=94450 $D=0
M960 246 242 240 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=89820 $D=0
M961 247 243 241 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=94450 $D=0
M962 8 246 716 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=89820 $D=0
M963 8 247 717 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=94450 $D=0
M964 248 716 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=89820 $D=0
M965 249 717 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=94450 $D=0
M966 246 16 248 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=89820 $D=0
M967 247 16 249 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=94450 $D=0
M968 248 244 250 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=89820 $D=0
M969 249 245 251 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=94450 $D=0
M970 254 252 248 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=89820 $D=0
M971 255 253 249 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=94450 $D=0
M972 252 18 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=89820 $D=0
M973 253 18 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=94450 $D=0
M974 8 19 256 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=89820 $D=0
M975 8 19 257 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=94450 $D=0
M976 258 20 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=89820 $D=0
M977 259 20 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=94450 $D=0
M978 260 256 240 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=89820 $D=0
M979 261 257 241 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=94450 $D=0
M980 8 260 718 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=89820 $D=0
M981 8 261 719 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=94450 $D=0
M982 262 718 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=89820 $D=0
M983 263 719 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=94450 $D=0
M984 260 19 262 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=89820 $D=0
M985 261 19 263 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=94450 $D=0
M986 262 258 250 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=89820 $D=0
M987 263 259 251 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=94450 $D=0
M988 254 264 262 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=89820 $D=0
M989 255 265 263 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=94450 $D=0
M990 264 21 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=89820 $D=0
M991 265 21 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=94450 $D=0
M992 8 22 266 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=89820 $D=0
M993 8 22 267 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=94450 $D=0
M994 268 23 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=89820 $D=0
M995 269 23 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=94450 $D=0
M996 270 266 240 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=89820 $D=0
M997 271 267 241 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=94450 $D=0
M998 8 270 720 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=89820 $D=0
M999 8 271 721 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=94450 $D=0
M1000 272 720 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=89820 $D=0
M1001 273 721 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=94450 $D=0
M1002 270 22 272 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=89820 $D=0
M1003 271 22 273 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=94450 $D=0
M1004 272 268 250 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=89820 $D=0
M1005 273 269 251 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=94450 $D=0
M1006 254 274 272 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=89820 $D=0
M1007 255 275 273 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=94450 $D=0
M1008 274 24 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=89820 $D=0
M1009 275 24 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=94450 $D=0
M1010 8 25 276 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=89820 $D=0
M1011 8 25 277 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=94450 $D=0
M1012 278 26 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=89820 $D=0
M1013 279 26 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=94450 $D=0
M1014 280 276 240 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=89820 $D=0
M1015 281 277 241 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=94450 $D=0
M1016 8 280 722 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=89820 $D=0
M1017 8 281 723 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=94450 $D=0
M1018 282 722 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=89820 $D=0
M1019 283 723 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=94450 $D=0
M1020 280 25 282 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=89820 $D=0
M1021 281 25 283 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=94450 $D=0
M1022 282 278 250 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=89820 $D=0
M1023 283 279 251 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=94450 $D=0
M1024 254 284 282 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=89820 $D=0
M1025 255 285 283 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=94450 $D=0
M1026 284 27 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=89820 $D=0
M1027 285 27 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=94450 $D=0
M1028 8 28 286 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=89820 $D=0
M1029 8 28 287 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=94450 $D=0
M1030 288 29 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=89820 $D=0
M1031 289 29 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=94450 $D=0
M1032 290 286 240 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=89820 $D=0
M1033 291 287 241 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=94450 $D=0
M1034 8 290 724 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=89820 $D=0
M1035 8 291 725 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=94450 $D=0
M1036 292 724 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=89820 $D=0
M1037 293 725 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=94450 $D=0
M1038 290 28 292 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=89820 $D=0
M1039 291 28 293 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=94450 $D=0
M1040 292 288 250 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=89820 $D=0
M1041 293 289 251 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=94450 $D=0
M1042 254 294 292 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=89820 $D=0
M1043 255 295 293 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=94450 $D=0
M1044 294 30 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=89820 $D=0
M1045 295 30 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=94450 $D=0
M1046 8 31 296 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=89820 $D=0
M1047 8 31 297 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=94450 $D=0
M1048 298 32 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=89820 $D=0
M1049 299 32 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=94450 $D=0
M1050 300 296 240 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=89820 $D=0
M1051 301 297 241 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=94450 $D=0
M1052 8 300 726 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=89820 $D=0
M1053 8 301 727 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=94450 $D=0
M1054 302 726 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=89820 $D=0
M1055 303 727 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=94450 $D=0
M1056 300 31 302 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=89820 $D=0
M1057 301 31 303 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=94450 $D=0
M1058 302 298 250 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=89820 $D=0
M1059 303 299 251 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=94450 $D=0
M1060 254 304 302 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=89820 $D=0
M1061 255 305 303 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=94450 $D=0
M1062 304 33 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=89820 $D=0
M1063 305 33 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=94450 $D=0
M1064 8 34 306 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=89820 $D=0
M1065 8 34 307 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=94450 $D=0
M1066 308 35 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=89820 $D=0
M1067 309 35 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=94450 $D=0
M1068 310 306 240 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=89820 $D=0
M1069 311 307 241 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=94450 $D=0
M1070 8 310 728 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=89820 $D=0
M1071 8 311 729 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=94450 $D=0
M1072 312 728 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=89820 $D=0
M1073 313 729 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=94450 $D=0
M1074 310 34 312 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=89820 $D=0
M1075 311 34 313 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=94450 $D=0
M1076 312 308 250 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=89820 $D=0
M1077 313 309 251 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=94450 $D=0
M1078 254 314 312 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=89820 $D=0
M1079 255 315 313 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=94450 $D=0
M1080 314 36 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=89820 $D=0
M1081 315 36 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=94450 $D=0
M1082 8 37 316 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=89820 $D=0
M1083 8 37 317 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=94450 $D=0
M1084 318 38 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=89820 $D=0
M1085 319 38 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=94450 $D=0
M1086 320 316 240 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=89820 $D=0
M1087 321 317 241 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=94450 $D=0
M1088 8 320 730 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=89820 $D=0
M1089 8 321 731 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=94450 $D=0
M1090 322 730 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=89820 $D=0
M1091 323 731 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=94450 $D=0
M1092 320 37 322 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=89820 $D=0
M1093 321 37 323 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=94450 $D=0
M1094 322 318 250 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=89820 $D=0
M1095 323 319 251 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=94450 $D=0
M1096 254 324 322 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=89820 $D=0
M1097 255 325 323 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=94450 $D=0
M1098 324 39 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=89820 $D=0
M1099 325 39 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=94450 $D=0
M1100 8 40 326 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=89820 $D=0
M1101 8 40 327 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=94450 $D=0
M1102 328 41 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=89820 $D=0
M1103 329 41 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=94450 $D=0
M1104 330 326 240 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=89820 $D=0
M1105 331 327 241 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=94450 $D=0
M1106 8 330 732 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=89820 $D=0
M1107 8 331 733 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=94450 $D=0
M1108 332 732 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=89820 $D=0
M1109 333 733 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=94450 $D=0
M1110 330 40 332 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=89820 $D=0
M1111 331 40 333 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=94450 $D=0
M1112 332 328 250 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=89820 $D=0
M1113 333 329 251 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=94450 $D=0
M1114 254 334 332 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=89820 $D=0
M1115 255 335 333 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=94450 $D=0
M1116 334 42 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=89820 $D=0
M1117 335 42 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=94450 $D=0
M1118 8 43 336 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=89820 $D=0
M1119 8 43 337 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=94450 $D=0
M1120 338 44 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=89820 $D=0
M1121 339 44 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=94450 $D=0
M1122 340 336 240 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=89820 $D=0
M1123 341 337 241 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=94450 $D=0
M1124 8 340 734 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=89820 $D=0
M1125 8 341 735 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=94450 $D=0
M1126 342 734 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=89820 $D=0
M1127 343 735 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=94450 $D=0
M1128 340 43 342 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=89820 $D=0
M1129 341 43 343 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=94450 $D=0
M1130 342 338 250 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=89820 $D=0
M1131 343 339 251 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=94450 $D=0
M1132 254 344 342 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=89820 $D=0
M1133 255 345 343 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=94450 $D=0
M1134 344 45 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=89820 $D=0
M1135 345 45 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=94450 $D=0
M1136 8 46 346 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=89820 $D=0
M1137 8 46 347 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=94450 $D=0
M1138 348 47 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=89820 $D=0
M1139 349 47 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=94450 $D=0
M1140 350 346 240 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=89820 $D=0
M1141 351 347 241 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=94450 $D=0
M1142 8 350 736 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=89820 $D=0
M1143 8 351 737 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=94450 $D=0
M1144 352 736 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=89820 $D=0
M1145 353 737 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=94450 $D=0
M1146 350 46 352 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=89820 $D=0
M1147 351 46 353 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=94450 $D=0
M1148 352 348 250 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=89820 $D=0
M1149 353 349 251 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=94450 $D=0
M1150 254 354 352 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=89820 $D=0
M1151 255 355 353 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=94450 $D=0
M1152 354 48 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=89820 $D=0
M1153 355 48 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=94450 $D=0
M1154 8 49 356 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=89820 $D=0
M1155 8 49 357 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=94450 $D=0
M1156 358 50 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=89820 $D=0
M1157 359 50 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=94450 $D=0
M1158 360 356 240 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=89820 $D=0
M1159 361 357 241 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=94450 $D=0
M1160 8 360 738 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=89820 $D=0
M1161 8 361 739 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=94450 $D=0
M1162 362 738 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=89820 $D=0
M1163 363 739 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=94450 $D=0
M1164 360 49 362 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=89820 $D=0
M1165 361 49 363 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=94450 $D=0
M1166 362 358 250 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=89820 $D=0
M1167 363 359 251 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=94450 $D=0
M1168 254 364 362 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=89820 $D=0
M1169 255 365 363 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=94450 $D=0
M1170 364 51 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=89820 $D=0
M1171 365 51 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=94450 $D=0
M1172 8 52 366 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=89820 $D=0
M1173 8 52 367 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=94450 $D=0
M1174 368 53 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=89820 $D=0
M1175 369 53 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=94450 $D=0
M1176 370 366 240 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=89820 $D=0
M1177 371 367 241 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=94450 $D=0
M1178 8 370 740 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=89820 $D=0
M1179 8 371 741 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=94450 $D=0
M1180 372 740 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=89820 $D=0
M1181 373 741 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=94450 $D=0
M1182 370 52 372 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=89820 $D=0
M1183 371 52 373 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=94450 $D=0
M1184 372 368 250 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=89820 $D=0
M1185 373 369 251 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=94450 $D=0
M1186 254 374 372 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=89820 $D=0
M1187 255 375 373 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=94450 $D=0
M1188 374 54 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=89820 $D=0
M1189 375 54 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=94450 $D=0
M1190 8 55 376 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=89820 $D=0
M1191 8 55 377 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=94450 $D=0
M1192 378 56 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=89820 $D=0
M1193 379 56 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=94450 $D=0
M1194 380 376 240 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=89820 $D=0
M1195 381 377 241 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=94450 $D=0
M1196 8 380 742 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=89820 $D=0
M1197 8 381 743 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=94450 $D=0
M1198 382 742 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=89820 $D=0
M1199 383 743 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=94450 $D=0
M1200 380 55 382 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=89820 $D=0
M1201 381 55 383 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=94450 $D=0
M1202 382 378 250 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=89820 $D=0
M1203 383 379 251 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=94450 $D=0
M1204 254 384 382 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=89820 $D=0
M1205 255 385 383 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=94450 $D=0
M1206 384 57 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=89820 $D=0
M1207 385 57 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=94450 $D=0
M1208 8 58 386 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=89820 $D=0
M1209 8 58 387 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=94450 $D=0
M1210 388 59 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=89820 $D=0
M1211 389 59 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=94450 $D=0
M1212 390 386 240 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=89820 $D=0
M1213 391 387 241 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=94450 $D=0
M1214 8 390 744 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=89820 $D=0
M1215 8 391 745 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=94450 $D=0
M1216 392 744 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=89820 $D=0
M1217 393 745 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=94450 $D=0
M1218 390 58 392 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=89820 $D=0
M1219 391 58 393 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=94450 $D=0
M1220 392 388 250 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=89820 $D=0
M1221 393 389 251 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=94450 $D=0
M1222 254 394 392 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=89820 $D=0
M1223 255 395 393 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=94450 $D=0
M1224 394 60 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=89820 $D=0
M1225 395 60 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=94450 $D=0
M1226 8 61 396 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=89820 $D=0
M1227 8 61 397 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=94450 $D=0
M1228 398 62 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=89820 $D=0
M1229 399 62 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=94450 $D=0
M1230 400 396 240 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=89820 $D=0
M1231 401 397 241 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=94450 $D=0
M1232 8 400 746 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=89820 $D=0
M1233 8 401 747 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=94450 $D=0
M1234 402 746 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=89820 $D=0
M1235 403 747 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=94450 $D=0
M1236 400 61 402 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=89820 $D=0
M1237 401 61 403 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=94450 $D=0
M1238 402 398 250 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=89820 $D=0
M1239 403 399 251 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=94450 $D=0
M1240 254 404 402 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=89820 $D=0
M1241 255 405 403 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=94450 $D=0
M1242 404 63 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=89820 $D=0
M1243 405 63 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=94450 $D=0
M1244 8 64 406 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=89820 $D=0
M1245 8 64 407 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=94450 $D=0
M1246 408 65 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=89820 $D=0
M1247 409 65 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=94450 $D=0
M1248 410 406 240 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=89820 $D=0
M1249 411 407 241 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=94450 $D=0
M1250 8 410 748 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=89820 $D=0
M1251 8 411 749 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=94450 $D=0
M1252 412 748 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=89820 $D=0
M1253 413 749 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=94450 $D=0
M1254 410 64 412 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=89820 $D=0
M1255 411 64 413 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=94450 $D=0
M1256 412 408 250 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=89820 $D=0
M1257 413 409 251 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=94450 $D=0
M1258 254 414 412 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=89820 $D=0
M1259 255 415 413 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=94450 $D=0
M1260 414 66 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=89820 $D=0
M1261 415 66 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=94450 $D=0
M1262 8 67 416 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=89820 $D=0
M1263 8 67 417 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=94450 $D=0
M1264 418 68 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=89820 $D=0
M1265 419 68 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=94450 $D=0
M1266 420 416 240 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=89820 $D=0
M1267 421 417 241 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=94450 $D=0
M1268 8 420 750 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=89820 $D=0
M1269 8 421 751 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=94450 $D=0
M1270 422 750 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=89820 $D=0
M1271 423 751 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=94450 $D=0
M1272 420 67 422 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=89820 $D=0
M1273 421 67 423 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=94450 $D=0
M1274 422 418 250 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=89820 $D=0
M1275 423 419 251 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=94450 $D=0
M1276 254 424 422 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=89820 $D=0
M1277 255 425 423 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=94450 $D=0
M1278 424 69 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=89820 $D=0
M1279 425 69 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=94450 $D=0
M1280 8 70 426 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=89820 $D=0
M1281 8 70 427 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=94450 $D=0
M1282 428 71 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=89820 $D=0
M1283 429 71 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=94450 $D=0
M1284 430 426 240 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=89820 $D=0
M1285 431 427 241 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=94450 $D=0
M1286 8 430 752 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=89820 $D=0
M1287 8 431 753 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=94450 $D=0
M1288 432 752 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=89820 $D=0
M1289 433 753 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=94450 $D=0
M1290 430 70 432 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=89820 $D=0
M1291 431 70 433 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=94450 $D=0
M1292 432 428 250 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=89820 $D=0
M1293 433 429 251 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=94450 $D=0
M1294 254 434 432 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=89820 $D=0
M1295 255 435 433 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=94450 $D=0
M1296 434 72 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=89820 $D=0
M1297 435 72 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=94450 $D=0
M1298 8 73 436 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=89820 $D=0
M1299 8 73 437 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=94450 $D=0
M1300 438 74 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=89820 $D=0
M1301 439 74 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=94450 $D=0
M1302 440 436 240 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=89820 $D=0
M1303 441 437 241 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=94450 $D=0
M1304 8 440 754 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=89820 $D=0
M1305 8 441 755 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=94450 $D=0
M1306 442 754 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=89820 $D=0
M1307 443 755 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=94450 $D=0
M1308 440 73 442 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=89820 $D=0
M1309 441 73 443 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=94450 $D=0
M1310 442 438 250 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=89820 $D=0
M1311 443 439 251 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=94450 $D=0
M1312 254 444 442 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=89820 $D=0
M1313 255 445 443 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=94450 $D=0
M1314 444 75 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=89820 $D=0
M1315 445 75 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=94450 $D=0
M1316 8 76 446 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=89820 $D=0
M1317 8 76 447 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=94450 $D=0
M1318 448 77 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=89820 $D=0
M1319 449 77 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=94450 $D=0
M1320 450 446 240 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=89820 $D=0
M1321 451 447 241 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=94450 $D=0
M1322 8 450 756 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=89820 $D=0
M1323 8 451 757 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=94450 $D=0
M1324 452 756 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=89820 $D=0
M1325 453 757 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=94450 $D=0
M1326 450 76 452 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=89820 $D=0
M1327 451 76 453 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=94450 $D=0
M1328 452 448 250 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=89820 $D=0
M1329 453 449 251 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=94450 $D=0
M1330 254 454 452 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=89820 $D=0
M1331 255 455 453 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=94450 $D=0
M1332 454 78 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=89820 $D=0
M1333 455 78 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=94450 $D=0
M1334 8 79 456 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=89820 $D=0
M1335 8 79 457 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=94450 $D=0
M1336 458 80 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=89820 $D=0
M1337 459 80 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=94450 $D=0
M1338 460 456 240 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=89820 $D=0
M1339 461 457 241 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=94450 $D=0
M1340 8 460 758 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=89820 $D=0
M1341 8 461 759 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=94450 $D=0
M1342 462 758 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=89820 $D=0
M1343 463 759 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=94450 $D=0
M1344 460 79 462 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=89820 $D=0
M1345 461 79 463 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=94450 $D=0
M1346 462 458 250 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=89820 $D=0
M1347 463 459 251 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=94450 $D=0
M1348 254 464 462 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=89820 $D=0
M1349 255 465 463 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=94450 $D=0
M1350 464 81 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=89820 $D=0
M1351 465 81 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=94450 $D=0
M1352 8 82 466 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=89820 $D=0
M1353 8 82 467 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=94450 $D=0
M1354 468 83 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=89820 $D=0
M1355 469 83 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=94450 $D=0
M1356 470 466 240 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=89820 $D=0
M1357 471 467 241 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=94450 $D=0
M1358 8 470 760 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=89820 $D=0
M1359 8 471 761 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=94450 $D=0
M1360 472 760 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=89820 $D=0
M1361 473 761 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=94450 $D=0
M1362 470 82 472 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=89820 $D=0
M1363 471 82 473 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=94450 $D=0
M1364 472 468 250 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=89820 $D=0
M1365 473 469 251 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=94450 $D=0
M1366 254 474 472 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=89820 $D=0
M1367 255 475 473 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=94450 $D=0
M1368 474 84 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=89820 $D=0
M1369 475 84 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=94450 $D=0
M1370 8 85 476 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=89820 $D=0
M1371 8 85 477 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=94450 $D=0
M1372 478 86 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=89820 $D=0
M1373 479 86 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=94450 $D=0
M1374 480 476 240 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=89820 $D=0
M1375 481 477 241 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=94450 $D=0
M1376 8 480 762 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=89820 $D=0
M1377 8 481 763 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=94450 $D=0
M1378 482 762 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=89820 $D=0
M1379 483 763 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=94450 $D=0
M1380 480 85 482 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=89820 $D=0
M1381 481 85 483 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=94450 $D=0
M1382 482 478 250 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=89820 $D=0
M1383 483 479 251 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=94450 $D=0
M1384 254 484 482 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=89820 $D=0
M1385 255 485 483 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=94450 $D=0
M1386 484 87 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=89820 $D=0
M1387 485 87 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=94450 $D=0
M1388 8 88 486 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=89820 $D=0
M1389 8 88 487 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=94450 $D=0
M1390 488 89 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=89820 $D=0
M1391 489 89 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=94450 $D=0
M1392 490 486 240 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=89820 $D=0
M1393 491 487 241 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=94450 $D=0
M1394 8 490 764 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=89820 $D=0
M1395 8 491 765 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=94450 $D=0
M1396 492 764 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=89820 $D=0
M1397 493 765 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=94450 $D=0
M1398 490 88 492 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=89820 $D=0
M1399 491 88 493 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=94450 $D=0
M1400 492 488 250 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=89820 $D=0
M1401 493 489 251 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=94450 $D=0
M1402 254 494 492 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=89820 $D=0
M1403 255 495 493 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=94450 $D=0
M1404 494 90 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=89820 $D=0
M1405 495 90 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=94450 $D=0
M1406 8 91 496 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=89820 $D=0
M1407 8 91 497 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=94450 $D=0
M1408 498 92 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=89820 $D=0
M1409 499 92 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=94450 $D=0
M1410 500 496 240 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=89820 $D=0
M1411 501 497 241 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=94450 $D=0
M1412 8 500 766 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=89820 $D=0
M1413 8 501 767 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=94450 $D=0
M1414 502 766 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=89820 $D=0
M1415 503 767 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=94450 $D=0
M1416 500 91 502 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=89820 $D=0
M1417 501 91 503 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=94450 $D=0
M1418 502 498 250 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=89820 $D=0
M1419 503 499 251 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=94450 $D=0
M1420 254 504 502 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=89820 $D=0
M1421 255 505 503 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=94450 $D=0
M1422 504 93 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=89820 $D=0
M1423 505 93 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=94450 $D=0
M1424 8 94 506 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=89820 $D=0
M1425 8 94 507 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=94450 $D=0
M1426 508 95 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=89820 $D=0
M1427 509 95 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=94450 $D=0
M1428 510 506 240 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=89820 $D=0
M1429 511 507 241 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=94450 $D=0
M1430 8 510 768 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=89820 $D=0
M1431 8 511 769 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=94450 $D=0
M1432 512 768 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=89820 $D=0
M1433 513 769 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=94450 $D=0
M1434 510 94 512 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=89820 $D=0
M1435 511 94 513 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=94450 $D=0
M1436 512 508 250 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=89820 $D=0
M1437 513 509 251 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=94450 $D=0
M1438 254 514 512 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=89820 $D=0
M1439 255 515 513 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=94450 $D=0
M1440 514 96 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=89820 $D=0
M1441 515 96 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=94450 $D=0
M1442 8 97 516 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=89820 $D=0
M1443 8 97 517 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=94450 $D=0
M1444 518 98 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=89820 $D=0
M1445 519 98 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=94450 $D=0
M1446 520 516 240 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=89820 $D=0
M1447 521 517 241 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=94450 $D=0
M1448 8 520 770 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=89820 $D=0
M1449 8 521 771 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=94450 $D=0
M1450 522 770 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=89820 $D=0
M1451 523 771 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=94450 $D=0
M1452 520 97 522 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=89820 $D=0
M1453 521 97 523 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=94450 $D=0
M1454 522 518 250 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=89820 $D=0
M1455 523 519 251 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=94450 $D=0
M1456 254 524 522 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=89820 $D=0
M1457 255 525 523 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=94450 $D=0
M1458 524 99 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=89820 $D=0
M1459 525 99 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=94450 $D=0
M1460 8 100 526 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=89820 $D=0
M1461 8 100 527 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=94450 $D=0
M1462 528 101 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=89820 $D=0
M1463 529 101 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=94450 $D=0
M1464 530 526 240 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=89820 $D=0
M1465 531 527 241 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=94450 $D=0
M1466 8 530 772 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=89820 $D=0
M1467 8 531 773 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=94450 $D=0
M1468 532 772 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=89820 $D=0
M1469 533 773 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=94450 $D=0
M1470 530 100 532 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=89820 $D=0
M1471 531 100 533 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=94450 $D=0
M1472 532 528 250 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=89820 $D=0
M1473 533 529 251 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=94450 $D=0
M1474 254 534 532 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=89820 $D=0
M1475 255 535 533 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=94450 $D=0
M1476 534 102 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=89820 $D=0
M1477 535 102 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=94450 $D=0
M1478 8 103 536 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=89820 $D=0
M1479 8 103 537 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=94450 $D=0
M1480 538 104 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=89820 $D=0
M1481 539 104 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=94450 $D=0
M1482 540 536 240 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=89820 $D=0
M1483 541 537 241 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=94450 $D=0
M1484 8 540 774 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=89820 $D=0
M1485 8 541 775 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=94450 $D=0
M1486 542 774 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=89820 $D=0
M1487 543 775 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=94450 $D=0
M1488 540 103 542 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=89820 $D=0
M1489 541 103 543 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=94450 $D=0
M1490 542 538 250 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=89820 $D=0
M1491 543 539 251 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=94450 $D=0
M1492 254 544 542 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=89820 $D=0
M1493 255 545 543 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=94450 $D=0
M1494 544 105 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=89820 $D=0
M1495 545 105 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=94450 $D=0
M1496 8 106 546 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=89820 $D=0
M1497 8 106 547 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=94450 $D=0
M1498 548 107 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=89820 $D=0
M1499 549 107 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=94450 $D=0
M1500 550 546 240 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=89820 $D=0
M1501 551 547 241 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=94450 $D=0
M1502 8 550 776 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=89820 $D=0
M1503 8 551 777 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=94450 $D=0
M1504 552 776 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=89820 $D=0
M1505 553 777 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=94450 $D=0
M1506 550 106 552 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=89820 $D=0
M1507 551 106 553 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=94450 $D=0
M1508 552 548 250 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=89820 $D=0
M1509 553 549 251 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=94450 $D=0
M1510 254 554 552 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=89820 $D=0
M1511 255 555 553 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=94450 $D=0
M1512 554 108 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=89820 $D=0
M1513 555 108 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=94450 $D=0
M1514 8 109 556 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=89820 $D=0
M1515 8 109 557 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=94450 $D=0
M1516 558 110 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=89820 $D=0
M1517 559 110 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=94450 $D=0
M1518 5 558 250 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=89820 $D=0
M1519 5 559 251 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=94450 $D=0
M1520 254 556 5 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=89820 $D=0
M1521 255 557 5 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=94450 $D=0
M1522 8 562 560 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=89820 $D=0
M1523 8 563 561 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=94450 $D=0
M1524 562 111 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=89820 $D=0
M1525 563 111 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=94450 $D=0
M1526 778 250 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=89820 $D=0
M1527 779 251 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=94450 $D=0
M1528 564 562 778 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=89820 $D=0
M1529 565 563 779 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=94450 $D=0
M1530 8 564 566 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=89820 $D=0
M1531 8 565 567 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=94450 $D=0
M1532 780 566 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=89820 $D=0
M1533 781 567 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=94450 $D=0
M1534 564 560 780 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=89820 $D=0
M1535 565 561 781 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=94450 $D=0
M1536 8 570 568 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=89820 $D=0
M1537 8 571 569 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=94450 $D=0
M1538 570 111 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=89820 $D=0
M1539 571 111 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=94450 $D=0
M1540 782 254 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=89820 $D=0
M1541 783 255 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=94450 $D=0
M1542 572 570 782 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=89820 $D=0
M1543 573 571 783 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=94450 $D=0
M1544 8 572 112 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=89820 $D=0
M1545 8 573 113 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=94450 $D=0
M1546 784 112 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=89820 $D=0
M1547 785 113 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=94450 $D=0
M1548 572 568 784 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=89820 $D=0
M1549 573 569 785 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=94450 $D=0
M1550 574 118 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=89820 $D=0
M1551 575 118 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=94450 $D=0
M1552 576 118 566 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=89820 $D=0
M1553 577 118 567 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=94450 $D=0
M1554 119 574 576 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=89820 $D=0
M1555 120 575 577 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=94450 $D=0
M1556 578 121 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=89820 $D=0
M1557 579 121 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=94450 $D=0
M1558 580 121 112 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=89820 $D=0
M1559 581 121 113 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=94450 $D=0
M1560 786 578 580 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=89820 $D=0
M1561 787 579 581 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=94450 $D=0
M1562 8 112 786 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=89820 $D=0
M1563 8 113 787 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=94450 $D=0
M1564 582 123 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=89820 $D=0
M1565 583 123 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=94450 $D=0
M1566 584 123 580 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=89820 $D=0
M1567 585 123 581 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=94450 $D=0
M1568 10 582 584 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=89820 $D=0
M1569 11 583 585 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=94450 $D=0
M1570 587 586 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=89820 $D=0
M1571 588 124 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=94450 $D=0
M1572 8 591 589 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=89820 $D=0
M1573 8 592 590 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=94450 $D=0
M1574 593 576 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=89820 $D=0
M1575 594 577 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=94450 $D=0
M1576 591 576 586 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=89820 $D=0
M1577 592 577 124 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=94450 $D=0
M1578 587 593 591 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=89820 $D=0
M1579 588 594 592 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=94450 $D=0
M1580 595 589 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=89820 $D=0
M1581 596 590 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=94450 $D=0
M1582 127 589 584 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=89820 $D=0
M1583 586 590 585 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=94450 $D=0
M1584 576 595 127 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=89820 $D=0
M1585 577 596 586 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=94450 $D=0
M1586 597 127 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=89820 $D=0
M1587 598 586 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=94450 $D=0
M1588 599 589 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=89820 $D=0
M1589 600 590 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=94450 $D=0
M1590 601 589 597 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=89820 $D=0
M1591 602 590 598 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=94450 $D=0
M1592 584 599 601 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=89820 $D=0
M1593 585 600 602 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=94450 $D=0
M1594 798 576 8 8 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=89460 $D=0
M1595 799 577 8 8 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=94090 $D=0
M1596 603 584 798 8 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=89460 $D=0
M1597 604 585 799 8 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=94090 $D=0
M1598 605 601 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=89820 $D=0
M1599 606 602 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=94450 $D=0
M1600 607 576 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=89820 $D=0
M1601 608 577 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=94450 $D=0
M1602 8 584 607 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=89820 $D=0
M1603 8 585 608 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=94450 $D=0
M1604 609 576 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=89820 $D=0
M1605 610 577 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=94450 $D=0
M1606 8 584 609 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=89820 $D=0
M1607 8 585 610 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=94450 $D=0
M1608 800 576 8 8 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=89640 $D=0
M1609 801 577 8 8 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=94270 $D=0
M1610 613 584 800 8 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=89640 $D=0
M1611 614 585 801 8 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=94270 $D=0
M1612 8 609 613 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=89820 $D=0
M1613 8 610 614 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=94450 $D=0
M1614 615 128 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=89820 $D=0
M1615 616 128 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=94450 $D=0
M1616 617 128 603 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=89820 $D=0
M1617 618 128 604 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=94450 $D=0
M1618 607 615 617 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=89820 $D=0
M1619 608 616 618 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=94450 $D=0
M1620 619 128 605 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=89820 $D=0
M1621 620 128 606 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=94450 $D=0
M1622 613 615 619 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=89820 $D=0
M1623 614 616 620 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=94450 $D=0
M1624 621 129 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=89820 $D=0
M1625 622 129 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=94450 $D=0
M1626 623 129 619 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=89820 $D=0
M1627 624 129 620 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=94450 $D=0
M1628 617 621 623 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=89820 $D=0
M1629 618 622 624 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=94450 $D=0
M1630 12 623 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=89820 $D=0
M1631 13 624 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=94450 $D=0
M1632 625 130 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=89820 $D=0
M1633 626 130 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=94450 $D=0
M1634 627 130 131 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=89820 $D=0
M1635 628 130 132 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=94450 $D=0
M1636 133 625 627 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=89820 $D=0
M1637 134 626 628 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=94450 $D=0
M1638 629 130 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=89820 $D=0
M1639 630 130 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=94450 $D=0
M1640 631 130 135 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=89820 $D=0
M1641 632 130 136 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=94450 $D=0
M1642 137 629 631 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=89820 $D=0
M1643 138 630 632 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=94450 $D=0
M1644 633 130 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=89820 $D=0
M1645 634 130 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=94450 $D=0
M1646 635 130 139 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=89820 $D=0
M1647 636 130 140 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=94450 $D=0
M1648 114 633 635 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=89820 $D=0
M1649 116 634 636 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=94450 $D=0
M1650 637 130 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=89820 $D=0
M1651 638 130 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=94450 $D=0
M1652 639 130 141 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=89820 $D=0
M1653 640 130 142 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=94450 $D=0
M1654 115 637 639 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=89820 $D=0
M1655 117 638 640 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=94450 $D=0
M1656 641 130 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=89820 $D=0
M1657 642 130 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=94450 $D=0
M1658 643 130 5 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=89820 $D=0
M1659 644 130 5 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=94450 $D=0
M1660 143 641 643 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=89820 $D=0
M1661 144 642 644 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=94450 $D=0
M1662 8 576 788 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=89820 $D=0
M1663 8 577 789 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=94450 $D=0
M1664 134 788 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=89820 $D=0
M1665 131 789 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=94450 $D=0
M1666 645 145 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=89820 $D=0
M1667 646 145 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=94450 $D=0
M1668 146 145 134 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=89820 $D=0
M1669 147 145 131 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=94450 $D=0
M1670 627 645 146 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=89820 $D=0
M1671 628 646 147 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=94450 $D=0
M1672 647 148 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=89820 $D=0
M1673 648 148 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=94450 $D=0
M1674 122 148 146 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=89820 $D=0
M1675 149 148 147 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=94450 $D=0
M1676 631 647 122 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=89820 $D=0
M1677 632 648 149 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=94450 $D=0
M1678 649 150 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=89820 $D=0
M1679 650 150 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=94450 $D=0
M1680 125 150 122 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=89820 $D=0
M1681 126 150 149 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=94450 $D=0
M1682 635 649 125 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=89820 $D=0
M1683 636 650 126 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=94450 $D=0
M1684 651 151 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=89820 $D=0
M1685 652 151 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=94450 $D=0
M1686 152 151 125 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=89820 $D=0
M1687 153 151 126 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=94450 $D=0
M1688 639 651 152 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=89820 $D=0
M1689 640 652 153 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=94450 $D=0
M1690 653 154 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=89820 $D=0
M1691 654 154 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=94450 $D=0
M1692 226 154 152 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=89820 $D=0
M1693 227 154 153 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=94450 $D=0
M1694 643 653 226 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=89820 $D=0
M1695 644 654 227 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=94450 $D=0
M1696 655 155 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=89820 $D=0
M1697 656 155 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=94450 $D=0
M1698 657 155 112 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=89820 $D=0
M1699 658 155 113 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=94450 $D=0
M1700 10 655 657 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=89820 $D=0
M1701 11 656 658 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=94450 $D=0
M1702 659 566 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=89820 $D=0
M1703 660 567 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=94450 $D=0
M1704 8 657 659 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=89820 $D=0
M1705 8 658 660 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=94450 $D=0
M1706 802 566 8 8 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=89640 $D=0
M1707 803 567 8 8 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=94270 $D=0
M1708 663 657 802 8 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=89640 $D=0
M1709 664 658 803 8 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=94270 $D=0
M1710 8 659 663 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=89820 $D=0
M1711 8 660 664 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=94450 $D=0
M1712 790 156 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=89820 $D=0
M1713 791 665 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=94450 $D=0
M1714 8 663 790 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=89820 $D=0
M1715 8 664 791 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=94450 $D=0
M1716 665 790 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=89820 $D=0
M1717 157 791 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=94450 $D=0
M1718 804 566 8 8 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=89460 $D=0
M1719 805 567 8 8 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=94090 $D=0
M1720 666 668 804 8 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=89460 $D=0
M1721 667 669 805 8 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=94090 $D=0
M1722 668 657 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=89820 $D=0
M1723 669 658 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=94450 $D=0
M1724 670 666 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=89820 $D=0
M1725 671 667 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=94450 $D=0
M1726 8 156 670 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=89820 $D=0
M1727 8 665 671 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=94450 $D=0
M1728 673 158 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=89820 $D=0
M1729 674 672 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=94450 $D=0
M1730 672 670 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=89820 $D=0
M1731 159 671 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=94450 $D=0
M1732 8 673 672 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=89820 $D=0
M1733 8 674 159 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=94450 $D=0
M1734 676 675 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=89820 $D=0
M1735 677 160 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=94450 $D=0
M1736 8 680 678 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=89820 $D=0
M1737 8 681 679 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=94450 $D=0
M1738 682 119 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=89820 $D=0
M1739 683 120 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=94450 $D=0
M1740 680 119 675 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=89820 $D=0
M1741 681 120 160 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=94450 $D=0
M1742 676 682 680 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=89820 $D=0
M1743 677 683 681 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=94450 $D=0
M1744 684 678 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=89820 $D=0
M1745 685 679 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=94450 $D=0
M1746 161 678 5 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=89820 $D=0
M1747 675 679 5 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=94450 $D=0
M1748 119 684 161 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=89820 $D=0
M1749 120 685 675 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=94450 $D=0
M1750 686 161 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=89820 $D=0
M1751 687 675 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=94450 $D=0
M1752 688 678 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=89820 $D=0
M1753 689 679 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=94450 $D=0
M1754 228 678 686 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=89820 $D=0
M1755 229 679 687 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=94450 $D=0
M1756 5 688 228 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=89820 $D=0
M1757 5 689 229 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=94450 $D=0
M1758 690 162 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=89820 $D=0
M1759 691 162 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=94450 $D=0
M1760 692 162 228 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=89820 $D=0
M1761 693 162 229 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=94450 $D=0
M1762 12 690 692 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=89820 $D=0
M1763 13 691 693 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=94450 $D=0
M1764 694 163 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=89820 $D=0
M1765 695 163 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=94450 $D=0
M1766 696 163 692 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=89820 $D=0
M1767 697 163 693 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=94450 $D=0
M1768 5 694 696 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=89820 $D=0
M1769 5 695 697 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=94450 $D=0
M1770 698 111 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=89820 $D=0
M1771 699 111 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=94450 $D=0
M1772 8 698 700 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=89820 $D=0
M1773 8 699 701 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=94450 $D=0
M1774 702 111 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=89820 $D=0
M1775 703 111 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=94450 $D=0
M1776 704 700 696 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=89820 $D=0
M1777 705 701 697 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=94450 $D=0
M1778 8 704 792 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=89820 $D=0
M1779 8 705 793 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=94450 $D=0
M1780 706 792 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=89820 $D=0
M1781 707 793 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=94450 $D=0
M1782 704 698 706 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=89820 $D=0
M1783 705 699 707 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=94450 $D=0
M1784 708 702 706 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=89820 $D=0
M1785 709 703 707 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=94450 $D=0
M1786 8 712 710 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=89820 $D=0
M1787 8 713 711 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=94450 $D=0
M1788 712 111 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=89820 $D=0
M1789 713 111 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=94450 $D=0
M1790 794 708 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=89820 $D=0
M1791 795 709 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=94450 $D=0
M1792 714 712 794 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=89820 $D=0
M1793 715 713 795 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=94450 $D=0
M1794 8 714 119 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=89820 $D=0
M1795 8 715 120 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=94450 $D=0
M1796 796 119 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=89820 $D=0
M1797 797 120 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=94450 $D=0
M1798 714 710 796 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=89820 $D=0
M1799 715 711 797 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=94450 $D=0
.ENDS
***************************************
.SUBCKT ICV_30 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163
** N=822 EP=163 IP=1514 FDC=1800
M0 206 1 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=79310 $D=1
M1 207 1 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=83940 $D=1
M2 208 206 2 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=79310 $D=1
M3 209 207 3 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=83940 $D=1
M4 5 1 208 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=79310 $D=1
M5 5 1 209 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=83940 $D=1
M6 210 206 4 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=79310 $D=1
M7 211 207 4 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=83940 $D=1
M8 2 1 210 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=79310 $D=1
M9 3 1 211 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=83940 $D=1
M10 212 206 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=79310 $D=1
M11 213 207 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=83940 $D=1
M12 2 1 212 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=79310 $D=1
M13 3 1 213 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=83940 $D=1
M14 216 214 212 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=79310 $D=1
M15 217 215 213 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=83940 $D=1
M16 214 6 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=79310 $D=1
M17 215 6 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=83940 $D=1
M18 218 214 210 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=79310 $D=1
M19 219 215 211 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=83940 $D=1
M20 208 6 218 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=79310 $D=1
M21 209 6 219 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=83940 $D=1
M22 220 7 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=79310 $D=1
M23 221 7 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=83940 $D=1
M24 222 220 218 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=79310 $D=1
M25 223 221 219 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=83940 $D=1
M26 216 7 222 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=79310 $D=1
M27 217 7 223 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=83940 $D=1
M28 224 9 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=79310 $D=1
M29 225 9 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=83940 $D=1
M30 226 224 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=79310 $D=1
M31 227 225 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=83940 $D=1
M32 10 9 226 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=79310 $D=1
M33 11 9 227 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=83940 $D=1
M34 228 224 12 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=79310 $D=1
M35 229 225 13 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=83940 $D=1
M36 230 9 228 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=79310 $D=1
M37 231 9 229 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=83940 $D=1
M38 234 224 232 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=79310 $D=1
M39 235 225 233 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=83940 $D=1
M40 222 9 234 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=79310 $D=1
M41 223 9 235 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=83940 $D=1
M42 238 236 234 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=79310 $D=1
M43 239 237 235 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=83940 $D=1
M44 236 14 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=79310 $D=1
M45 237 14 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=83940 $D=1
M46 240 236 228 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=79310 $D=1
M47 241 237 229 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=83940 $D=1
M48 226 14 240 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=79310 $D=1
M49 227 14 241 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=83940 $D=1
M50 242 15 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=79310 $D=1
M51 243 15 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=83940 $D=1
M52 244 242 240 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=79310 $D=1
M53 245 243 241 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=83940 $D=1
M54 238 15 244 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=79310 $D=1
M55 239 15 245 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=83940 $D=1
M56 5 16 246 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=79310 $D=1
M57 5 16 247 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=83940 $D=1
M58 248 17 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=79310 $D=1
M59 249 17 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=83940 $D=1
M60 250 16 244 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=79310 $D=1
M61 251 16 245 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=83940 $D=1
M62 5 250 721 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=79310 $D=1
M63 5 251 722 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=83940 $D=1
M64 252 721 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=79310 $D=1
M65 253 722 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=83940 $D=1
M66 250 246 252 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=79310 $D=1
M67 251 247 253 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=83940 $D=1
M68 252 17 254 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=79310 $D=1
M69 253 17 255 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=83940 $D=1
M70 258 18 252 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=79310 $D=1
M71 259 18 253 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=83940 $D=1
M72 256 18 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=79310 $D=1
M73 257 18 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=83940 $D=1
M74 5 19 260 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=79310 $D=1
M75 5 19 261 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=83940 $D=1
M76 262 20 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=79310 $D=1
M77 263 20 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=83940 $D=1
M78 264 19 244 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=79310 $D=1
M79 265 19 245 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=83940 $D=1
M80 5 264 723 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=79310 $D=1
M81 5 265 724 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=83940 $D=1
M82 266 723 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=79310 $D=1
M83 267 724 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=83940 $D=1
M84 264 260 266 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=79310 $D=1
M85 265 261 267 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=83940 $D=1
M86 266 20 254 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=79310 $D=1
M87 267 20 255 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=83940 $D=1
M88 258 21 266 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=79310 $D=1
M89 259 21 267 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=83940 $D=1
M90 268 21 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=79310 $D=1
M91 269 21 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=83940 $D=1
M92 5 22 270 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=79310 $D=1
M93 5 22 271 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=83940 $D=1
M94 272 23 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=79310 $D=1
M95 273 23 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=83940 $D=1
M96 274 22 244 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=79310 $D=1
M97 275 22 245 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=83940 $D=1
M98 5 274 725 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=79310 $D=1
M99 5 275 726 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=83940 $D=1
M100 276 725 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=79310 $D=1
M101 277 726 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=83940 $D=1
M102 274 270 276 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=79310 $D=1
M103 275 271 277 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=83940 $D=1
M104 276 23 254 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=79310 $D=1
M105 277 23 255 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=83940 $D=1
M106 258 24 276 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=79310 $D=1
M107 259 24 277 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=83940 $D=1
M108 278 24 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=79310 $D=1
M109 279 24 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=83940 $D=1
M110 5 25 280 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=79310 $D=1
M111 5 25 281 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=83940 $D=1
M112 282 26 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=79310 $D=1
M113 283 26 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=83940 $D=1
M114 284 25 244 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=79310 $D=1
M115 285 25 245 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=83940 $D=1
M116 5 284 727 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=79310 $D=1
M117 5 285 728 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=83940 $D=1
M118 286 727 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=79310 $D=1
M119 287 728 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=83940 $D=1
M120 284 280 286 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=79310 $D=1
M121 285 281 287 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=83940 $D=1
M122 286 26 254 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=79310 $D=1
M123 287 26 255 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=83940 $D=1
M124 258 27 286 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=79310 $D=1
M125 259 27 287 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=83940 $D=1
M126 288 27 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=79310 $D=1
M127 289 27 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=83940 $D=1
M128 5 28 290 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=79310 $D=1
M129 5 28 291 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=83940 $D=1
M130 292 29 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=79310 $D=1
M131 293 29 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=83940 $D=1
M132 294 28 244 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=79310 $D=1
M133 295 28 245 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=83940 $D=1
M134 5 294 729 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=79310 $D=1
M135 5 295 730 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=83940 $D=1
M136 296 729 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=79310 $D=1
M137 297 730 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=83940 $D=1
M138 294 290 296 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=79310 $D=1
M139 295 291 297 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=83940 $D=1
M140 296 29 254 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=79310 $D=1
M141 297 29 255 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=83940 $D=1
M142 258 30 296 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=79310 $D=1
M143 259 30 297 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=83940 $D=1
M144 298 30 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=79310 $D=1
M145 299 30 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=83940 $D=1
M146 5 31 300 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=79310 $D=1
M147 5 31 301 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=83940 $D=1
M148 302 32 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=79310 $D=1
M149 303 32 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=83940 $D=1
M150 304 31 244 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=79310 $D=1
M151 305 31 245 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=83940 $D=1
M152 5 304 731 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=79310 $D=1
M153 5 305 732 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=83940 $D=1
M154 306 731 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=79310 $D=1
M155 307 732 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=83940 $D=1
M156 304 300 306 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=79310 $D=1
M157 305 301 307 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=83940 $D=1
M158 306 32 254 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=79310 $D=1
M159 307 32 255 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=83940 $D=1
M160 258 33 306 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=79310 $D=1
M161 259 33 307 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=83940 $D=1
M162 308 33 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=79310 $D=1
M163 309 33 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=83940 $D=1
M164 5 34 310 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=79310 $D=1
M165 5 34 311 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=83940 $D=1
M166 312 35 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=79310 $D=1
M167 313 35 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=83940 $D=1
M168 314 34 244 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=79310 $D=1
M169 315 34 245 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=83940 $D=1
M170 5 314 733 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=79310 $D=1
M171 5 315 734 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=83940 $D=1
M172 316 733 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=79310 $D=1
M173 317 734 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=83940 $D=1
M174 314 310 316 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=79310 $D=1
M175 315 311 317 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=83940 $D=1
M176 316 35 254 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=79310 $D=1
M177 317 35 255 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=83940 $D=1
M178 258 36 316 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=79310 $D=1
M179 259 36 317 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=83940 $D=1
M180 318 36 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=79310 $D=1
M181 319 36 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=83940 $D=1
M182 5 37 320 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=79310 $D=1
M183 5 37 321 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=83940 $D=1
M184 322 38 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=79310 $D=1
M185 323 38 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=83940 $D=1
M186 324 37 244 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=79310 $D=1
M187 325 37 245 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=83940 $D=1
M188 5 324 735 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=79310 $D=1
M189 5 325 736 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=83940 $D=1
M190 326 735 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=79310 $D=1
M191 327 736 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=83940 $D=1
M192 324 320 326 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=79310 $D=1
M193 325 321 327 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=83940 $D=1
M194 326 38 254 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=79310 $D=1
M195 327 38 255 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=83940 $D=1
M196 258 39 326 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=79310 $D=1
M197 259 39 327 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=83940 $D=1
M198 328 39 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=79310 $D=1
M199 329 39 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=83940 $D=1
M200 5 40 330 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=79310 $D=1
M201 5 40 331 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=83940 $D=1
M202 332 41 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=79310 $D=1
M203 333 41 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=83940 $D=1
M204 334 40 244 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=79310 $D=1
M205 335 40 245 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=83940 $D=1
M206 5 334 737 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=79310 $D=1
M207 5 335 738 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=83940 $D=1
M208 336 737 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=79310 $D=1
M209 337 738 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=83940 $D=1
M210 334 330 336 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=79310 $D=1
M211 335 331 337 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=83940 $D=1
M212 336 41 254 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=79310 $D=1
M213 337 41 255 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=83940 $D=1
M214 258 42 336 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=79310 $D=1
M215 259 42 337 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=83940 $D=1
M216 338 42 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=79310 $D=1
M217 339 42 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=83940 $D=1
M218 5 43 340 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=79310 $D=1
M219 5 43 341 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=83940 $D=1
M220 342 44 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=79310 $D=1
M221 343 44 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=83940 $D=1
M222 344 43 244 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=79310 $D=1
M223 345 43 245 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=83940 $D=1
M224 5 344 739 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=79310 $D=1
M225 5 345 740 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=83940 $D=1
M226 346 739 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=79310 $D=1
M227 347 740 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=83940 $D=1
M228 344 340 346 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=79310 $D=1
M229 345 341 347 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=83940 $D=1
M230 346 44 254 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=79310 $D=1
M231 347 44 255 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=83940 $D=1
M232 258 45 346 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=79310 $D=1
M233 259 45 347 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=83940 $D=1
M234 348 45 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=79310 $D=1
M235 349 45 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=83940 $D=1
M236 5 46 350 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=79310 $D=1
M237 5 46 351 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=83940 $D=1
M238 352 47 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=79310 $D=1
M239 353 47 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=83940 $D=1
M240 354 46 244 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=79310 $D=1
M241 355 46 245 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=83940 $D=1
M242 5 354 741 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=79310 $D=1
M243 5 355 742 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=83940 $D=1
M244 356 741 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=79310 $D=1
M245 357 742 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=83940 $D=1
M246 354 350 356 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=79310 $D=1
M247 355 351 357 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=83940 $D=1
M248 356 47 254 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=79310 $D=1
M249 357 47 255 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=83940 $D=1
M250 258 48 356 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=79310 $D=1
M251 259 48 357 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=83940 $D=1
M252 358 48 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=79310 $D=1
M253 359 48 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=83940 $D=1
M254 5 49 360 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=79310 $D=1
M255 5 49 361 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=83940 $D=1
M256 362 50 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=79310 $D=1
M257 363 50 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=83940 $D=1
M258 364 49 244 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=79310 $D=1
M259 365 49 245 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=83940 $D=1
M260 5 364 743 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=79310 $D=1
M261 5 365 744 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=83940 $D=1
M262 366 743 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=79310 $D=1
M263 367 744 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=83940 $D=1
M264 364 360 366 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=79310 $D=1
M265 365 361 367 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=83940 $D=1
M266 366 50 254 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=79310 $D=1
M267 367 50 255 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=83940 $D=1
M268 258 51 366 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=79310 $D=1
M269 259 51 367 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=83940 $D=1
M270 368 51 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=79310 $D=1
M271 369 51 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=83940 $D=1
M272 5 52 370 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=79310 $D=1
M273 5 52 371 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=83940 $D=1
M274 372 53 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=79310 $D=1
M275 373 53 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=83940 $D=1
M276 374 52 244 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=79310 $D=1
M277 375 52 245 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=83940 $D=1
M278 5 374 745 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=79310 $D=1
M279 5 375 746 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=83940 $D=1
M280 376 745 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=79310 $D=1
M281 377 746 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=83940 $D=1
M282 374 370 376 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=79310 $D=1
M283 375 371 377 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=83940 $D=1
M284 376 53 254 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=79310 $D=1
M285 377 53 255 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=83940 $D=1
M286 258 54 376 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=79310 $D=1
M287 259 54 377 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=83940 $D=1
M288 378 54 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=79310 $D=1
M289 379 54 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=83940 $D=1
M290 5 55 380 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=79310 $D=1
M291 5 55 381 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=83940 $D=1
M292 382 56 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=79310 $D=1
M293 383 56 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=83940 $D=1
M294 384 55 244 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=79310 $D=1
M295 385 55 245 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=83940 $D=1
M296 5 384 747 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=79310 $D=1
M297 5 385 748 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=83940 $D=1
M298 386 747 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=79310 $D=1
M299 387 748 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=83940 $D=1
M300 384 380 386 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=79310 $D=1
M301 385 381 387 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=83940 $D=1
M302 386 56 254 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=79310 $D=1
M303 387 56 255 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=83940 $D=1
M304 258 57 386 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=79310 $D=1
M305 259 57 387 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=83940 $D=1
M306 388 57 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=79310 $D=1
M307 389 57 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=83940 $D=1
M308 5 58 390 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=79310 $D=1
M309 5 58 391 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=83940 $D=1
M310 392 59 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=79310 $D=1
M311 393 59 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=83940 $D=1
M312 394 58 244 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=79310 $D=1
M313 395 58 245 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=83940 $D=1
M314 5 394 749 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=79310 $D=1
M315 5 395 750 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=83940 $D=1
M316 396 749 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=79310 $D=1
M317 397 750 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=83940 $D=1
M318 394 390 396 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=79310 $D=1
M319 395 391 397 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=83940 $D=1
M320 396 59 254 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=79310 $D=1
M321 397 59 255 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=83940 $D=1
M322 258 60 396 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=79310 $D=1
M323 259 60 397 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=83940 $D=1
M324 398 60 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=79310 $D=1
M325 399 60 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=83940 $D=1
M326 5 61 400 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=79310 $D=1
M327 5 61 401 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=83940 $D=1
M328 402 62 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=79310 $D=1
M329 403 62 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=83940 $D=1
M330 404 61 244 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=79310 $D=1
M331 405 61 245 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=83940 $D=1
M332 5 404 751 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=79310 $D=1
M333 5 405 752 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=83940 $D=1
M334 406 751 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=79310 $D=1
M335 407 752 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=83940 $D=1
M336 404 400 406 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=79310 $D=1
M337 405 401 407 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=83940 $D=1
M338 406 62 254 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=79310 $D=1
M339 407 62 255 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=83940 $D=1
M340 258 63 406 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=79310 $D=1
M341 259 63 407 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=83940 $D=1
M342 408 63 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=79310 $D=1
M343 409 63 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=83940 $D=1
M344 5 64 410 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=79310 $D=1
M345 5 64 411 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=83940 $D=1
M346 412 65 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=79310 $D=1
M347 413 65 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=83940 $D=1
M348 414 64 244 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=79310 $D=1
M349 415 64 245 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=83940 $D=1
M350 5 414 753 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=79310 $D=1
M351 5 415 754 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=83940 $D=1
M352 416 753 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=79310 $D=1
M353 417 754 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=83940 $D=1
M354 414 410 416 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=79310 $D=1
M355 415 411 417 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=83940 $D=1
M356 416 65 254 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=79310 $D=1
M357 417 65 255 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=83940 $D=1
M358 258 66 416 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=79310 $D=1
M359 259 66 417 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=83940 $D=1
M360 418 66 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=79310 $D=1
M361 419 66 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=83940 $D=1
M362 5 67 420 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=79310 $D=1
M363 5 67 421 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=83940 $D=1
M364 422 68 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=79310 $D=1
M365 423 68 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=83940 $D=1
M366 424 67 244 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=79310 $D=1
M367 425 67 245 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=83940 $D=1
M368 5 424 755 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=79310 $D=1
M369 5 425 756 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=83940 $D=1
M370 426 755 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=79310 $D=1
M371 427 756 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=83940 $D=1
M372 424 420 426 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=79310 $D=1
M373 425 421 427 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=83940 $D=1
M374 426 68 254 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=79310 $D=1
M375 427 68 255 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=83940 $D=1
M376 258 69 426 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=79310 $D=1
M377 259 69 427 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=83940 $D=1
M378 428 69 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=79310 $D=1
M379 429 69 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=83940 $D=1
M380 5 70 430 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=79310 $D=1
M381 5 70 431 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=83940 $D=1
M382 432 71 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=79310 $D=1
M383 433 71 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=83940 $D=1
M384 434 70 244 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=79310 $D=1
M385 435 70 245 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=83940 $D=1
M386 5 434 757 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=79310 $D=1
M387 5 435 758 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=83940 $D=1
M388 436 757 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=79310 $D=1
M389 437 758 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=83940 $D=1
M390 434 430 436 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=79310 $D=1
M391 435 431 437 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=83940 $D=1
M392 436 71 254 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=79310 $D=1
M393 437 71 255 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=83940 $D=1
M394 258 72 436 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=79310 $D=1
M395 259 72 437 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=83940 $D=1
M396 438 72 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=79310 $D=1
M397 439 72 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=83940 $D=1
M398 5 73 440 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=79310 $D=1
M399 5 73 441 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=83940 $D=1
M400 442 74 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=79310 $D=1
M401 443 74 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=83940 $D=1
M402 444 73 244 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=79310 $D=1
M403 445 73 245 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=83940 $D=1
M404 5 444 759 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=79310 $D=1
M405 5 445 760 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=83940 $D=1
M406 446 759 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=79310 $D=1
M407 447 760 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=83940 $D=1
M408 444 440 446 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=79310 $D=1
M409 445 441 447 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=83940 $D=1
M410 446 74 254 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=79310 $D=1
M411 447 74 255 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=83940 $D=1
M412 258 75 446 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=79310 $D=1
M413 259 75 447 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=83940 $D=1
M414 448 75 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=79310 $D=1
M415 449 75 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=83940 $D=1
M416 5 76 450 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=79310 $D=1
M417 5 76 451 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=83940 $D=1
M418 452 77 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=79310 $D=1
M419 453 77 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=83940 $D=1
M420 454 76 244 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=79310 $D=1
M421 455 76 245 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=83940 $D=1
M422 5 454 761 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=79310 $D=1
M423 5 455 762 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=83940 $D=1
M424 456 761 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=79310 $D=1
M425 457 762 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=83940 $D=1
M426 454 450 456 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=79310 $D=1
M427 455 451 457 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=83940 $D=1
M428 456 77 254 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=79310 $D=1
M429 457 77 255 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=83940 $D=1
M430 258 78 456 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=79310 $D=1
M431 259 78 457 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=83940 $D=1
M432 458 78 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=79310 $D=1
M433 459 78 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=83940 $D=1
M434 5 79 460 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=79310 $D=1
M435 5 79 461 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=83940 $D=1
M436 462 80 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=79310 $D=1
M437 463 80 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=83940 $D=1
M438 464 79 244 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=79310 $D=1
M439 465 79 245 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=83940 $D=1
M440 5 464 763 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=79310 $D=1
M441 5 465 764 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=83940 $D=1
M442 466 763 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=79310 $D=1
M443 467 764 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=83940 $D=1
M444 464 460 466 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=79310 $D=1
M445 465 461 467 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=83940 $D=1
M446 466 80 254 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=79310 $D=1
M447 467 80 255 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=83940 $D=1
M448 258 81 466 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=79310 $D=1
M449 259 81 467 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=83940 $D=1
M450 468 81 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=79310 $D=1
M451 469 81 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=83940 $D=1
M452 5 82 470 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=79310 $D=1
M453 5 82 471 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=83940 $D=1
M454 472 83 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=79310 $D=1
M455 473 83 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=83940 $D=1
M456 474 82 244 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=79310 $D=1
M457 475 82 245 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=83940 $D=1
M458 5 474 765 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=79310 $D=1
M459 5 475 766 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=83940 $D=1
M460 476 765 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=79310 $D=1
M461 477 766 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=83940 $D=1
M462 474 470 476 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=79310 $D=1
M463 475 471 477 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=83940 $D=1
M464 476 83 254 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=79310 $D=1
M465 477 83 255 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=83940 $D=1
M466 258 84 476 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=79310 $D=1
M467 259 84 477 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=83940 $D=1
M468 478 84 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=79310 $D=1
M469 479 84 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=83940 $D=1
M470 5 85 480 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=79310 $D=1
M471 5 85 481 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=83940 $D=1
M472 482 86 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=79310 $D=1
M473 483 86 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=83940 $D=1
M474 484 85 244 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=79310 $D=1
M475 485 85 245 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=83940 $D=1
M476 5 484 767 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=79310 $D=1
M477 5 485 768 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=83940 $D=1
M478 486 767 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=79310 $D=1
M479 487 768 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=83940 $D=1
M480 484 480 486 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=79310 $D=1
M481 485 481 487 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=83940 $D=1
M482 486 86 254 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=79310 $D=1
M483 487 86 255 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=83940 $D=1
M484 258 87 486 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=79310 $D=1
M485 259 87 487 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=83940 $D=1
M486 488 87 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=79310 $D=1
M487 489 87 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=83940 $D=1
M488 5 88 490 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=79310 $D=1
M489 5 88 491 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=83940 $D=1
M490 492 89 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=79310 $D=1
M491 493 89 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=83940 $D=1
M492 494 88 244 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=79310 $D=1
M493 495 88 245 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=83940 $D=1
M494 5 494 769 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=79310 $D=1
M495 5 495 770 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=83940 $D=1
M496 496 769 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=79310 $D=1
M497 497 770 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=83940 $D=1
M498 494 490 496 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=79310 $D=1
M499 495 491 497 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=83940 $D=1
M500 496 89 254 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=79310 $D=1
M501 497 89 255 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=83940 $D=1
M502 258 90 496 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=79310 $D=1
M503 259 90 497 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=83940 $D=1
M504 498 90 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=79310 $D=1
M505 499 90 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=83940 $D=1
M506 5 91 500 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=79310 $D=1
M507 5 91 501 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=83940 $D=1
M508 502 92 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=79310 $D=1
M509 503 92 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=83940 $D=1
M510 504 91 244 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=79310 $D=1
M511 505 91 245 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=83940 $D=1
M512 5 504 771 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=79310 $D=1
M513 5 505 772 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=83940 $D=1
M514 506 771 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=79310 $D=1
M515 507 772 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=83940 $D=1
M516 504 500 506 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=79310 $D=1
M517 505 501 507 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=83940 $D=1
M518 506 92 254 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=79310 $D=1
M519 507 92 255 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=83940 $D=1
M520 258 93 506 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=79310 $D=1
M521 259 93 507 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=83940 $D=1
M522 508 93 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=79310 $D=1
M523 509 93 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=83940 $D=1
M524 5 94 510 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=79310 $D=1
M525 5 94 511 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=83940 $D=1
M526 512 95 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=79310 $D=1
M527 513 95 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=83940 $D=1
M528 514 94 244 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=79310 $D=1
M529 515 94 245 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=83940 $D=1
M530 5 514 773 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=79310 $D=1
M531 5 515 774 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=83940 $D=1
M532 516 773 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=79310 $D=1
M533 517 774 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=83940 $D=1
M534 514 510 516 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=79310 $D=1
M535 515 511 517 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=83940 $D=1
M536 516 95 254 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=79310 $D=1
M537 517 95 255 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=83940 $D=1
M538 258 96 516 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=79310 $D=1
M539 259 96 517 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=83940 $D=1
M540 518 96 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=79310 $D=1
M541 519 96 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=83940 $D=1
M542 5 97 520 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=79310 $D=1
M543 5 97 521 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=83940 $D=1
M544 522 98 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=79310 $D=1
M545 523 98 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=83940 $D=1
M546 524 97 244 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=79310 $D=1
M547 525 97 245 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=83940 $D=1
M548 5 524 775 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=79310 $D=1
M549 5 525 776 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=83940 $D=1
M550 526 775 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=79310 $D=1
M551 527 776 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=83940 $D=1
M552 524 520 526 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=79310 $D=1
M553 525 521 527 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=83940 $D=1
M554 526 98 254 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=79310 $D=1
M555 527 98 255 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=83940 $D=1
M556 258 99 526 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=79310 $D=1
M557 259 99 527 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=83940 $D=1
M558 528 99 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=79310 $D=1
M559 529 99 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=83940 $D=1
M560 5 100 530 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=79310 $D=1
M561 5 100 531 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=83940 $D=1
M562 532 101 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=79310 $D=1
M563 533 101 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=83940 $D=1
M564 534 100 244 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=79310 $D=1
M565 535 100 245 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=83940 $D=1
M566 5 534 777 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=79310 $D=1
M567 5 535 778 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=83940 $D=1
M568 536 777 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=79310 $D=1
M569 537 778 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=83940 $D=1
M570 534 530 536 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=79310 $D=1
M571 535 531 537 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=83940 $D=1
M572 536 101 254 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=79310 $D=1
M573 537 101 255 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=83940 $D=1
M574 258 102 536 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=79310 $D=1
M575 259 102 537 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=83940 $D=1
M576 538 102 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=79310 $D=1
M577 539 102 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=83940 $D=1
M578 5 103 540 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=79310 $D=1
M579 5 103 541 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=83940 $D=1
M580 542 104 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=79310 $D=1
M581 543 104 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=83940 $D=1
M582 544 103 244 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=79310 $D=1
M583 545 103 245 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=83940 $D=1
M584 5 544 779 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=79310 $D=1
M585 5 545 780 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=83940 $D=1
M586 546 779 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=79310 $D=1
M587 547 780 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=83940 $D=1
M588 544 540 546 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=79310 $D=1
M589 545 541 547 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=83940 $D=1
M590 546 104 254 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=79310 $D=1
M591 547 104 255 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=83940 $D=1
M592 258 105 546 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=79310 $D=1
M593 259 105 547 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=83940 $D=1
M594 548 105 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=79310 $D=1
M595 549 105 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=83940 $D=1
M596 5 106 550 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=79310 $D=1
M597 5 106 551 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=83940 $D=1
M598 552 107 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=79310 $D=1
M599 553 107 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=83940 $D=1
M600 554 106 244 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=79310 $D=1
M601 555 106 245 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=83940 $D=1
M602 5 554 781 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=79310 $D=1
M603 5 555 782 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=83940 $D=1
M604 556 781 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=79310 $D=1
M605 557 782 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=83940 $D=1
M606 554 550 556 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=79310 $D=1
M607 555 551 557 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=83940 $D=1
M608 556 107 254 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=79310 $D=1
M609 557 107 255 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=83940 $D=1
M610 258 108 556 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=79310 $D=1
M611 259 108 557 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=83940 $D=1
M612 558 108 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=79310 $D=1
M613 559 108 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=83940 $D=1
M614 5 109 560 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=79310 $D=1
M615 5 109 561 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=83940 $D=1
M616 562 110 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=79310 $D=1
M617 563 110 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=83940 $D=1
M618 5 110 254 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=79310 $D=1
M619 5 110 255 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=83940 $D=1
M620 258 109 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=79310 $D=1
M621 259 109 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=83940 $D=1
M622 5 566 564 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=79310 $D=1
M623 5 567 565 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=83940 $D=1
M624 566 111 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=79310 $D=1
M625 567 111 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=83940 $D=1
M626 783 254 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=79310 $D=1
M627 784 255 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=83940 $D=1
M628 568 564 783 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=79310 $D=1
M629 569 565 784 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=83940 $D=1
M630 5 568 570 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=79310 $D=1
M631 5 569 571 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=83940 $D=1
M632 785 570 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=79310 $D=1
M633 786 571 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=83940 $D=1
M634 568 566 785 5 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=79310 $D=1
M635 569 567 786 5 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=83940 $D=1
M636 5 575 573 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=79310 $D=1
M637 5 576 574 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=83940 $D=1
M638 575 111 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=79310 $D=1
M639 576 111 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=83940 $D=1
M640 787 258 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=79310 $D=1
M641 788 259 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=83940 $D=1
M642 577 573 787 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=79310 $D=1
M643 578 574 788 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=83940 $D=1
M644 5 577 117 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=79310 $D=1
M645 5 578 118 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=83940 $D=1
M646 789 117 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=79310 $D=1
M647 790 118 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=83940 $D=1
M648 577 575 789 5 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=79310 $D=1
M649 578 576 790 5 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=83940 $D=1
M650 579 119 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=79310 $D=1
M651 580 119 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=83940 $D=1
M652 581 579 570 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=79310 $D=1
M653 582 580 571 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=83940 $D=1
M654 121 119 581 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=79310 $D=1
M655 122 119 582 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=83940 $D=1
M656 583 123 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=79310 $D=1
M657 584 123 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=83940 $D=1
M658 585 583 117 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=79310 $D=1
M659 586 584 118 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=83940 $D=1
M660 791 123 585 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=79310 $D=1
M661 792 123 586 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=83940 $D=1
M662 5 117 791 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=79310 $D=1
M663 5 118 792 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=83940 $D=1
M664 587 125 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=79310 $D=1
M665 588 125 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=83940 $D=1
M666 589 587 585 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=79310 $D=1
M667 590 588 586 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=83940 $D=1
M668 10 125 589 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=79310 $D=1
M669 11 125 590 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=83940 $D=1
M670 592 591 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=79310 $D=1
M671 593 126 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=83940 $D=1
M672 5 596 594 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=79310 $D=1
M673 5 597 595 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=83940 $D=1
M674 598 581 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=79310 $D=1
M675 599 582 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=83940 $D=1
M676 596 598 591 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=79310 $D=1
M677 597 599 126 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=83940 $D=1
M678 592 581 596 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=79310 $D=1
M679 593 582 597 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=83940 $D=1
M680 600 594 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=79310 $D=1
M681 601 595 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=83940 $D=1
M682 128 600 589 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=79310 $D=1
M683 591 601 590 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=83940 $D=1
M684 581 594 128 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=79310 $D=1
M685 582 595 591 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=83940 $D=1
M686 602 128 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=79310 $D=1
M687 603 591 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=83940 $D=1
M688 604 594 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=79310 $D=1
M689 605 595 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=83940 $D=1
M690 606 604 602 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=79310 $D=1
M691 607 605 603 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=83940 $D=1
M692 589 594 606 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=79310 $D=1
M693 590 595 607 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=83940 $D=1
M694 608 581 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=79310 $D=1
M695 609 582 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=83940 $D=1
M696 5 589 608 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=79310 $D=1
M697 5 590 609 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=83940 $D=1
M698 610 606 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=79310 $D=1
M699 611 607 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=83940 $D=1
M700 811 581 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=79310 $D=1
M701 812 582 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=83940 $D=1
M702 612 589 811 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=79310 $D=1
M703 613 590 812 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=83940 $D=1
M704 813 581 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=79310 $D=1
M705 814 582 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=83940 $D=1
M706 614 589 813 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=79310 $D=1
M707 615 590 814 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=83940 $D=1
M708 618 581 616 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=79310 $D=1
M709 619 582 617 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=83940 $D=1
M710 616 589 618 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=79310 $D=1
M711 617 590 619 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=83940 $D=1
M712 5 614 616 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=79310 $D=1
M713 5 615 617 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=83940 $D=1
M714 620 129 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=79310 $D=1
M715 621 129 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=83940 $D=1
M716 622 620 608 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=79310 $D=1
M717 623 621 609 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=83940 $D=1
M718 612 129 622 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=79310 $D=1
M719 613 129 623 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=83940 $D=1
M720 624 620 610 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=79310 $D=1
M721 625 621 611 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=83940 $D=1
M722 618 129 624 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=79310 $D=1
M723 619 129 625 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=83940 $D=1
M724 626 130 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=79310 $D=1
M725 627 130 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=83940 $D=1
M726 628 626 624 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=79310 $D=1
M727 629 627 625 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=83940 $D=1
M728 622 130 628 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=79310 $D=1
M729 623 130 629 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=83940 $D=1
M730 12 628 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=79310 $D=1
M731 13 629 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=83940 $D=1
M732 630 131 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=79310 $D=1
M733 631 131 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=83940 $D=1
M734 632 630 132 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=79310 $D=1
M735 633 631 133 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=83940 $D=1
M736 134 131 632 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=79310 $D=1
M737 135 131 633 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=83940 $D=1
M738 634 131 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=79310 $D=1
M739 635 131 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=83940 $D=1
M740 636 634 136 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=79310 $D=1
M741 637 635 137 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=83940 $D=1
M742 138 131 636 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=79310 $D=1
M743 139 131 637 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=83940 $D=1
M744 638 131 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=79310 $D=1
M745 639 131 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=83940 $D=1
M746 640 638 140 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=79310 $D=1
M747 641 639 141 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=83940 $D=1
M748 113 131 640 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=79310 $D=1
M749 115 131 641 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=83940 $D=1
M750 642 131 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=79310 $D=1
M751 643 131 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=83940 $D=1
M752 644 642 142 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=79310 $D=1
M753 645 643 143 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=83940 $D=1
M754 114 131 644 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=79310 $D=1
M755 116 131 645 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=83940 $D=1
M756 646 131 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=79310 $D=1
M757 647 131 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=83940 $D=1
M758 648 646 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=79310 $D=1
M759 649 647 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=83940 $D=1
M760 144 131 648 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=79310 $D=1
M761 145 131 649 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=83940 $D=1
M762 5 581 793 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=79310 $D=1
M763 5 582 794 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=83940 $D=1
M764 135 793 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=79310 $D=1
M765 132 794 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=83940 $D=1
M766 650 146 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=79310 $D=1
M767 651 146 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=83940 $D=1
M768 147 650 135 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=79310 $D=1
M769 148 651 132 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=83940 $D=1
M770 632 146 147 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=79310 $D=1
M771 633 146 148 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=83940 $D=1
M772 652 149 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=79310 $D=1
M773 653 149 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=83940 $D=1
M774 120 652 147 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=79310 $D=1
M775 124 653 148 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=83940 $D=1
M776 636 149 120 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=79310 $D=1
M777 637 149 124 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=83940 $D=1
M778 654 150 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=79310 $D=1
M779 655 150 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=83940 $D=1
M780 112 654 120 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=79310 $D=1
M781 127 655 124 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=83940 $D=1
M782 640 150 112 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=79310 $D=1
M783 641 150 127 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=83940 $D=1
M784 656 151 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=79310 $D=1
M785 657 151 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=83940 $D=1
M786 152 656 112 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=79310 $D=1
M787 153 657 127 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=83940 $D=1
M788 644 151 152 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=79310 $D=1
M789 645 151 153 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=83940 $D=1
M790 658 154 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=79310 $D=1
M791 659 154 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=83940 $D=1
M792 230 658 152 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=79310 $D=1
M793 231 659 153 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=83940 $D=1
M794 648 154 230 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=79310 $D=1
M795 649 154 231 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=83940 $D=1
M796 660 155 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=79310 $D=1
M797 661 155 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=83940 $D=1
M798 662 660 117 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=79310 $D=1
M799 663 661 118 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=83940 $D=1
M800 10 155 662 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=79310 $D=1
M801 11 155 663 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=83940 $D=1
M802 815 570 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=79310 $D=1
M803 816 571 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=83940 $D=1
M804 664 662 815 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=79310 $D=1
M805 665 663 816 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=83940 $D=1
M806 668 570 666 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=79310 $D=1
M807 669 571 667 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=83940 $D=1
M808 666 662 668 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=79310 $D=1
M809 667 663 669 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=83940 $D=1
M810 5 664 666 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=79310 $D=1
M811 5 665 667 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=83940 $D=1
M812 817 156 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=79310 $D=1
M813 818 670 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=83940 $D=1
M814 795 668 817 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=79310 $D=1
M815 796 669 818 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=83940 $D=1
M816 670 795 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=79310 $D=1
M817 157 796 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=83940 $D=1
M818 671 570 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=79310 $D=1
M819 672 571 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=83940 $D=1
M820 5 673 671 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=79310 $D=1
M821 5 674 672 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=83940 $D=1
M822 673 662 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=79310 $D=1
M823 674 663 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=83940 $D=1
M824 819 671 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=79310 $D=1
M825 820 672 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=83940 $D=1
M826 675 156 819 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=79310 $D=1
M827 676 670 820 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=83940 $D=1
M828 678 158 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=79310 $D=1
M829 679 677 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=83940 $D=1
M830 821 675 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=79310 $D=1
M831 822 676 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=83940 $D=1
M832 677 678 821 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=79310 $D=1
M833 159 679 822 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=83940 $D=1
M834 681 680 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=79310 $D=1
M835 682 160 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=83940 $D=1
M836 5 685 683 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=79310 $D=1
M837 5 686 684 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=83940 $D=1
M838 687 121 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=79310 $D=1
M839 688 122 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=83940 $D=1
M840 685 687 680 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=79310 $D=1
M841 686 688 160 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=83940 $D=1
M842 681 121 685 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=79310 $D=1
M843 682 122 686 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=83940 $D=1
M844 689 683 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=79310 $D=1
M845 690 684 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=83940 $D=1
M846 161 689 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=79310 $D=1
M847 680 690 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=83940 $D=1
M848 121 683 161 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=79310 $D=1
M849 122 684 680 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=83940 $D=1
M850 691 161 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=79310 $D=1
M851 692 680 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=83940 $D=1
M852 693 683 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=79310 $D=1
M853 694 684 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=83940 $D=1
M854 232 693 691 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=79310 $D=1
M855 233 694 692 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=83940 $D=1
M856 5 683 232 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=79310 $D=1
M857 5 684 233 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=83940 $D=1
M858 695 162 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=79310 $D=1
M859 696 162 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=83940 $D=1
M860 697 695 232 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=79310 $D=1
M861 698 696 233 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=83940 $D=1
M862 12 162 697 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=79310 $D=1
M863 13 162 698 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=83940 $D=1
M864 699 163 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=79310 $D=1
M865 700 163 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=83940 $D=1
M866 701 699 697 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=79310 $D=1
M867 702 700 698 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=83940 $D=1
M868 5 163 701 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=79310 $D=1
M869 5 163 702 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=83940 $D=1
M870 703 111 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=79310 $D=1
M871 704 111 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=83940 $D=1
M872 5 703 705 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=79310 $D=1
M873 5 704 706 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=83940 $D=1
M874 707 111 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=79310 $D=1
M875 708 111 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=83940 $D=1
M876 709 703 701 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=79310 $D=1
M877 710 704 702 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=83940 $D=1
M878 5 709 797 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=79310 $D=1
M879 5 710 798 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=83940 $D=1
M880 711 797 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=79310 $D=1
M881 712 798 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=83940 $D=1
M882 709 705 711 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=79310 $D=1
M883 710 706 712 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=83940 $D=1
M884 713 111 711 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=79310 $D=1
M885 714 111 712 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=83940 $D=1
M886 5 717 715 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=79310 $D=1
M887 5 718 716 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=83940 $D=1
M888 717 111 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=79310 $D=1
M889 718 111 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=83940 $D=1
M890 799 713 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=79310 $D=1
M891 800 714 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=83940 $D=1
M892 719 715 799 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=79310 $D=1
M893 720 716 800 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=83940 $D=1
M894 5 719 121 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=79310 $D=1
M895 5 720 122 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=83940 $D=1
M896 801 121 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=79310 $D=1
M897 802 122 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=83940 $D=1
M898 719 717 801 5 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=79310 $D=1
M899 720 718 802 5 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=83940 $D=1
M900 206 1 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=80560 $D=0
M901 207 1 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=85190 $D=0
M902 208 1 2 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=80560 $D=0
M903 209 1 3 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=85190 $D=0
M904 5 206 208 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=80560 $D=0
M905 5 207 209 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=85190 $D=0
M906 210 1 4 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=80560 $D=0
M907 211 1 4 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=85190 $D=0
M908 2 206 210 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=80560 $D=0
M909 3 207 211 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=85190 $D=0
M910 212 1 5 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=80560 $D=0
M911 213 1 5 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=85190 $D=0
M912 2 206 212 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=80560 $D=0
M913 3 207 213 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=85190 $D=0
M914 216 6 212 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=80560 $D=0
M915 217 6 213 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=85190 $D=0
M916 214 6 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=80560 $D=0
M917 215 6 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=85190 $D=0
M918 218 6 210 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=80560 $D=0
M919 219 6 211 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=85190 $D=0
M920 208 214 218 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=80560 $D=0
M921 209 215 219 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=85190 $D=0
M922 220 7 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=80560 $D=0
M923 221 7 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=85190 $D=0
M924 222 7 218 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=80560 $D=0
M925 223 7 219 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=85190 $D=0
M926 216 220 222 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=80560 $D=0
M927 217 221 223 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=85190 $D=0
M928 224 9 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=80560 $D=0
M929 225 9 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=85190 $D=0
M930 226 9 5 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=80560 $D=0
M931 227 9 5 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=85190 $D=0
M932 10 224 226 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=80560 $D=0
M933 11 225 227 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=85190 $D=0
M934 228 9 12 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=80560 $D=0
M935 229 9 13 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=85190 $D=0
M936 230 224 228 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=80560 $D=0
M937 231 225 229 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=85190 $D=0
M938 234 9 232 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=80560 $D=0
M939 235 9 233 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=85190 $D=0
M940 222 224 234 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=80560 $D=0
M941 223 225 235 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=85190 $D=0
M942 238 14 234 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=80560 $D=0
M943 239 14 235 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=85190 $D=0
M944 236 14 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=80560 $D=0
M945 237 14 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=85190 $D=0
M946 240 14 228 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=80560 $D=0
M947 241 14 229 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=85190 $D=0
M948 226 236 240 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=80560 $D=0
M949 227 237 241 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=85190 $D=0
M950 242 15 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=80560 $D=0
M951 243 15 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=85190 $D=0
M952 244 15 240 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=80560 $D=0
M953 245 15 241 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=85190 $D=0
M954 238 242 244 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=80560 $D=0
M955 239 243 245 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=85190 $D=0
M956 8 16 246 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=80560 $D=0
M957 8 16 247 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=85190 $D=0
M958 248 17 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=80560 $D=0
M959 249 17 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=85190 $D=0
M960 250 246 244 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=80560 $D=0
M961 251 247 245 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=85190 $D=0
M962 8 250 721 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=80560 $D=0
M963 8 251 722 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=85190 $D=0
M964 252 721 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=80560 $D=0
M965 253 722 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=85190 $D=0
M966 250 16 252 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=80560 $D=0
M967 251 16 253 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=85190 $D=0
M968 252 248 254 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=80560 $D=0
M969 253 249 255 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=85190 $D=0
M970 258 256 252 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=80560 $D=0
M971 259 257 253 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=85190 $D=0
M972 256 18 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=80560 $D=0
M973 257 18 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=85190 $D=0
M974 8 19 260 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=80560 $D=0
M975 8 19 261 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=85190 $D=0
M976 262 20 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=80560 $D=0
M977 263 20 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=85190 $D=0
M978 264 260 244 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=80560 $D=0
M979 265 261 245 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=85190 $D=0
M980 8 264 723 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=80560 $D=0
M981 8 265 724 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=85190 $D=0
M982 266 723 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=80560 $D=0
M983 267 724 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=85190 $D=0
M984 264 19 266 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=80560 $D=0
M985 265 19 267 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=85190 $D=0
M986 266 262 254 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=80560 $D=0
M987 267 263 255 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=85190 $D=0
M988 258 268 266 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=80560 $D=0
M989 259 269 267 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=85190 $D=0
M990 268 21 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=80560 $D=0
M991 269 21 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=85190 $D=0
M992 8 22 270 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=80560 $D=0
M993 8 22 271 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=85190 $D=0
M994 272 23 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=80560 $D=0
M995 273 23 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=85190 $D=0
M996 274 270 244 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=80560 $D=0
M997 275 271 245 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=85190 $D=0
M998 8 274 725 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=80560 $D=0
M999 8 275 726 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=85190 $D=0
M1000 276 725 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=80560 $D=0
M1001 277 726 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=85190 $D=0
M1002 274 22 276 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=80560 $D=0
M1003 275 22 277 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=85190 $D=0
M1004 276 272 254 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=80560 $D=0
M1005 277 273 255 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=85190 $D=0
M1006 258 278 276 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=80560 $D=0
M1007 259 279 277 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=85190 $D=0
M1008 278 24 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=80560 $D=0
M1009 279 24 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=85190 $D=0
M1010 8 25 280 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=80560 $D=0
M1011 8 25 281 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=85190 $D=0
M1012 282 26 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=80560 $D=0
M1013 283 26 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=85190 $D=0
M1014 284 280 244 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=80560 $D=0
M1015 285 281 245 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=85190 $D=0
M1016 8 284 727 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=80560 $D=0
M1017 8 285 728 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=85190 $D=0
M1018 286 727 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=80560 $D=0
M1019 287 728 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=85190 $D=0
M1020 284 25 286 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=80560 $D=0
M1021 285 25 287 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=85190 $D=0
M1022 286 282 254 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=80560 $D=0
M1023 287 283 255 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=85190 $D=0
M1024 258 288 286 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=80560 $D=0
M1025 259 289 287 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=85190 $D=0
M1026 288 27 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=80560 $D=0
M1027 289 27 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=85190 $D=0
M1028 8 28 290 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=80560 $D=0
M1029 8 28 291 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=85190 $D=0
M1030 292 29 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=80560 $D=0
M1031 293 29 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=85190 $D=0
M1032 294 290 244 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=80560 $D=0
M1033 295 291 245 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=85190 $D=0
M1034 8 294 729 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=80560 $D=0
M1035 8 295 730 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=85190 $D=0
M1036 296 729 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=80560 $D=0
M1037 297 730 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=85190 $D=0
M1038 294 28 296 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=80560 $D=0
M1039 295 28 297 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=85190 $D=0
M1040 296 292 254 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=80560 $D=0
M1041 297 293 255 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=85190 $D=0
M1042 258 298 296 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=80560 $D=0
M1043 259 299 297 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=85190 $D=0
M1044 298 30 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=80560 $D=0
M1045 299 30 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=85190 $D=0
M1046 8 31 300 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=80560 $D=0
M1047 8 31 301 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=85190 $D=0
M1048 302 32 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=80560 $D=0
M1049 303 32 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=85190 $D=0
M1050 304 300 244 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=80560 $D=0
M1051 305 301 245 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=85190 $D=0
M1052 8 304 731 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=80560 $D=0
M1053 8 305 732 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=85190 $D=0
M1054 306 731 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=80560 $D=0
M1055 307 732 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=85190 $D=0
M1056 304 31 306 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=80560 $D=0
M1057 305 31 307 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=85190 $D=0
M1058 306 302 254 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=80560 $D=0
M1059 307 303 255 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=85190 $D=0
M1060 258 308 306 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=80560 $D=0
M1061 259 309 307 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=85190 $D=0
M1062 308 33 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=80560 $D=0
M1063 309 33 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=85190 $D=0
M1064 8 34 310 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=80560 $D=0
M1065 8 34 311 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=85190 $D=0
M1066 312 35 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=80560 $D=0
M1067 313 35 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=85190 $D=0
M1068 314 310 244 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=80560 $D=0
M1069 315 311 245 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=85190 $D=0
M1070 8 314 733 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=80560 $D=0
M1071 8 315 734 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=85190 $D=0
M1072 316 733 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=80560 $D=0
M1073 317 734 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=85190 $D=0
M1074 314 34 316 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=80560 $D=0
M1075 315 34 317 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=85190 $D=0
M1076 316 312 254 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=80560 $D=0
M1077 317 313 255 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=85190 $D=0
M1078 258 318 316 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=80560 $D=0
M1079 259 319 317 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=85190 $D=0
M1080 318 36 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=80560 $D=0
M1081 319 36 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=85190 $D=0
M1082 8 37 320 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=80560 $D=0
M1083 8 37 321 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=85190 $D=0
M1084 322 38 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=80560 $D=0
M1085 323 38 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=85190 $D=0
M1086 324 320 244 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=80560 $D=0
M1087 325 321 245 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=85190 $D=0
M1088 8 324 735 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=80560 $D=0
M1089 8 325 736 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=85190 $D=0
M1090 326 735 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=80560 $D=0
M1091 327 736 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=85190 $D=0
M1092 324 37 326 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=80560 $D=0
M1093 325 37 327 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=85190 $D=0
M1094 326 322 254 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=80560 $D=0
M1095 327 323 255 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=85190 $D=0
M1096 258 328 326 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=80560 $D=0
M1097 259 329 327 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=85190 $D=0
M1098 328 39 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=80560 $D=0
M1099 329 39 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=85190 $D=0
M1100 8 40 330 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=80560 $D=0
M1101 8 40 331 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=85190 $D=0
M1102 332 41 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=80560 $D=0
M1103 333 41 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=85190 $D=0
M1104 334 330 244 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=80560 $D=0
M1105 335 331 245 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=85190 $D=0
M1106 8 334 737 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=80560 $D=0
M1107 8 335 738 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=85190 $D=0
M1108 336 737 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=80560 $D=0
M1109 337 738 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=85190 $D=0
M1110 334 40 336 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=80560 $D=0
M1111 335 40 337 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=85190 $D=0
M1112 336 332 254 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=80560 $D=0
M1113 337 333 255 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=85190 $D=0
M1114 258 338 336 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=80560 $D=0
M1115 259 339 337 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=85190 $D=0
M1116 338 42 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=80560 $D=0
M1117 339 42 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=85190 $D=0
M1118 8 43 340 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=80560 $D=0
M1119 8 43 341 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=85190 $D=0
M1120 342 44 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=80560 $D=0
M1121 343 44 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=85190 $D=0
M1122 344 340 244 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=80560 $D=0
M1123 345 341 245 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=85190 $D=0
M1124 8 344 739 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=80560 $D=0
M1125 8 345 740 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=85190 $D=0
M1126 346 739 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=80560 $D=0
M1127 347 740 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=85190 $D=0
M1128 344 43 346 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=80560 $D=0
M1129 345 43 347 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=85190 $D=0
M1130 346 342 254 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=80560 $D=0
M1131 347 343 255 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=85190 $D=0
M1132 258 348 346 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=80560 $D=0
M1133 259 349 347 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=85190 $D=0
M1134 348 45 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=80560 $D=0
M1135 349 45 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=85190 $D=0
M1136 8 46 350 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=80560 $D=0
M1137 8 46 351 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=85190 $D=0
M1138 352 47 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=80560 $D=0
M1139 353 47 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=85190 $D=0
M1140 354 350 244 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=80560 $D=0
M1141 355 351 245 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=85190 $D=0
M1142 8 354 741 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=80560 $D=0
M1143 8 355 742 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=85190 $D=0
M1144 356 741 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=80560 $D=0
M1145 357 742 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=85190 $D=0
M1146 354 46 356 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=80560 $D=0
M1147 355 46 357 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=85190 $D=0
M1148 356 352 254 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=80560 $D=0
M1149 357 353 255 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=85190 $D=0
M1150 258 358 356 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=80560 $D=0
M1151 259 359 357 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=85190 $D=0
M1152 358 48 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=80560 $D=0
M1153 359 48 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=85190 $D=0
M1154 8 49 360 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=80560 $D=0
M1155 8 49 361 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=85190 $D=0
M1156 362 50 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=80560 $D=0
M1157 363 50 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=85190 $D=0
M1158 364 360 244 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=80560 $D=0
M1159 365 361 245 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=85190 $D=0
M1160 8 364 743 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=80560 $D=0
M1161 8 365 744 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=85190 $D=0
M1162 366 743 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=80560 $D=0
M1163 367 744 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=85190 $D=0
M1164 364 49 366 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=80560 $D=0
M1165 365 49 367 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=85190 $D=0
M1166 366 362 254 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=80560 $D=0
M1167 367 363 255 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=85190 $D=0
M1168 258 368 366 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=80560 $D=0
M1169 259 369 367 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=85190 $D=0
M1170 368 51 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=80560 $D=0
M1171 369 51 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=85190 $D=0
M1172 8 52 370 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=80560 $D=0
M1173 8 52 371 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=85190 $D=0
M1174 372 53 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=80560 $D=0
M1175 373 53 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=85190 $D=0
M1176 374 370 244 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=80560 $D=0
M1177 375 371 245 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=85190 $D=0
M1178 8 374 745 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=80560 $D=0
M1179 8 375 746 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=85190 $D=0
M1180 376 745 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=80560 $D=0
M1181 377 746 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=85190 $D=0
M1182 374 52 376 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=80560 $D=0
M1183 375 52 377 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=85190 $D=0
M1184 376 372 254 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=80560 $D=0
M1185 377 373 255 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=85190 $D=0
M1186 258 378 376 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=80560 $D=0
M1187 259 379 377 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=85190 $D=0
M1188 378 54 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=80560 $D=0
M1189 379 54 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=85190 $D=0
M1190 8 55 380 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=80560 $D=0
M1191 8 55 381 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=85190 $D=0
M1192 382 56 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=80560 $D=0
M1193 383 56 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=85190 $D=0
M1194 384 380 244 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=80560 $D=0
M1195 385 381 245 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=85190 $D=0
M1196 8 384 747 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=80560 $D=0
M1197 8 385 748 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=85190 $D=0
M1198 386 747 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=80560 $D=0
M1199 387 748 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=85190 $D=0
M1200 384 55 386 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=80560 $D=0
M1201 385 55 387 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=85190 $D=0
M1202 386 382 254 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=80560 $D=0
M1203 387 383 255 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=85190 $D=0
M1204 258 388 386 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=80560 $D=0
M1205 259 389 387 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=85190 $D=0
M1206 388 57 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=80560 $D=0
M1207 389 57 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=85190 $D=0
M1208 8 58 390 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=80560 $D=0
M1209 8 58 391 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=85190 $D=0
M1210 392 59 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=80560 $D=0
M1211 393 59 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=85190 $D=0
M1212 394 390 244 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=80560 $D=0
M1213 395 391 245 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=85190 $D=0
M1214 8 394 749 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=80560 $D=0
M1215 8 395 750 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=85190 $D=0
M1216 396 749 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=80560 $D=0
M1217 397 750 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=85190 $D=0
M1218 394 58 396 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=80560 $D=0
M1219 395 58 397 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=85190 $D=0
M1220 396 392 254 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=80560 $D=0
M1221 397 393 255 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=85190 $D=0
M1222 258 398 396 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=80560 $D=0
M1223 259 399 397 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=85190 $D=0
M1224 398 60 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=80560 $D=0
M1225 399 60 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=85190 $D=0
M1226 8 61 400 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=80560 $D=0
M1227 8 61 401 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=85190 $D=0
M1228 402 62 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=80560 $D=0
M1229 403 62 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=85190 $D=0
M1230 404 400 244 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=80560 $D=0
M1231 405 401 245 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=85190 $D=0
M1232 8 404 751 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=80560 $D=0
M1233 8 405 752 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=85190 $D=0
M1234 406 751 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=80560 $D=0
M1235 407 752 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=85190 $D=0
M1236 404 61 406 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=80560 $D=0
M1237 405 61 407 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=85190 $D=0
M1238 406 402 254 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=80560 $D=0
M1239 407 403 255 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=85190 $D=0
M1240 258 408 406 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=80560 $D=0
M1241 259 409 407 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=85190 $D=0
M1242 408 63 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=80560 $D=0
M1243 409 63 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=85190 $D=0
M1244 8 64 410 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=80560 $D=0
M1245 8 64 411 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=85190 $D=0
M1246 412 65 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=80560 $D=0
M1247 413 65 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=85190 $D=0
M1248 414 410 244 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=80560 $D=0
M1249 415 411 245 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=85190 $D=0
M1250 8 414 753 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=80560 $D=0
M1251 8 415 754 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=85190 $D=0
M1252 416 753 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=80560 $D=0
M1253 417 754 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=85190 $D=0
M1254 414 64 416 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=80560 $D=0
M1255 415 64 417 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=85190 $D=0
M1256 416 412 254 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=80560 $D=0
M1257 417 413 255 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=85190 $D=0
M1258 258 418 416 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=80560 $D=0
M1259 259 419 417 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=85190 $D=0
M1260 418 66 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=80560 $D=0
M1261 419 66 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=85190 $D=0
M1262 8 67 420 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=80560 $D=0
M1263 8 67 421 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=85190 $D=0
M1264 422 68 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=80560 $D=0
M1265 423 68 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=85190 $D=0
M1266 424 420 244 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=80560 $D=0
M1267 425 421 245 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=85190 $D=0
M1268 8 424 755 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=80560 $D=0
M1269 8 425 756 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=85190 $D=0
M1270 426 755 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=80560 $D=0
M1271 427 756 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=85190 $D=0
M1272 424 67 426 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=80560 $D=0
M1273 425 67 427 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=85190 $D=0
M1274 426 422 254 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=80560 $D=0
M1275 427 423 255 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=85190 $D=0
M1276 258 428 426 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=80560 $D=0
M1277 259 429 427 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=85190 $D=0
M1278 428 69 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=80560 $D=0
M1279 429 69 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=85190 $D=0
M1280 8 70 430 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=80560 $D=0
M1281 8 70 431 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=85190 $D=0
M1282 432 71 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=80560 $D=0
M1283 433 71 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=85190 $D=0
M1284 434 430 244 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=80560 $D=0
M1285 435 431 245 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=85190 $D=0
M1286 8 434 757 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=80560 $D=0
M1287 8 435 758 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=85190 $D=0
M1288 436 757 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=80560 $D=0
M1289 437 758 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=85190 $D=0
M1290 434 70 436 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=80560 $D=0
M1291 435 70 437 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=85190 $D=0
M1292 436 432 254 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=80560 $D=0
M1293 437 433 255 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=85190 $D=0
M1294 258 438 436 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=80560 $D=0
M1295 259 439 437 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=85190 $D=0
M1296 438 72 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=80560 $D=0
M1297 439 72 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=85190 $D=0
M1298 8 73 440 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=80560 $D=0
M1299 8 73 441 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=85190 $D=0
M1300 442 74 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=80560 $D=0
M1301 443 74 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=85190 $D=0
M1302 444 440 244 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=80560 $D=0
M1303 445 441 245 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=85190 $D=0
M1304 8 444 759 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=80560 $D=0
M1305 8 445 760 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=85190 $D=0
M1306 446 759 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=80560 $D=0
M1307 447 760 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=85190 $D=0
M1308 444 73 446 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=80560 $D=0
M1309 445 73 447 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=85190 $D=0
M1310 446 442 254 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=80560 $D=0
M1311 447 443 255 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=85190 $D=0
M1312 258 448 446 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=80560 $D=0
M1313 259 449 447 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=85190 $D=0
M1314 448 75 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=80560 $D=0
M1315 449 75 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=85190 $D=0
M1316 8 76 450 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=80560 $D=0
M1317 8 76 451 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=85190 $D=0
M1318 452 77 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=80560 $D=0
M1319 453 77 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=85190 $D=0
M1320 454 450 244 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=80560 $D=0
M1321 455 451 245 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=85190 $D=0
M1322 8 454 761 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=80560 $D=0
M1323 8 455 762 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=85190 $D=0
M1324 456 761 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=80560 $D=0
M1325 457 762 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=85190 $D=0
M1326 454 76 456 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=80560 $D=0
M1327 455 76 457 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=85190 $D=0
M1328 456 452 254 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=80560 $D=0
M1329 457 453 255 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=85190 $D=0
M1330 258 458 456 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=80560 $D=0
M1331 259 459 457 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=85190 $D=0
M1332 458 78 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=80560 $D=0
M1333 459 78 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=85190 $D=0
M1334 8 79 460 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=80560 $D=0
M1335 8 79 461 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=85190 $D=0
M1336 462 80 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=80560 $D=0
M1337 463 80 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=85190 $D=0
M1338 464 460 244 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=80560 $D=0
M1339 465 461 245 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=85190 $D=0
M1340 8 464 763 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=80560 $D=0
M1341 8 465 764 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=85190 $D=0
M1342 466 763 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=80560 $D=0
M1343 467 764 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=85190 $D=0
M1344 464 79 466 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=80560 $D=0
M1345 465 79 467 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=85190 $D=0
M1346 466 462 254 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=80560 $D=0
M1347 467 463 255 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=85190 $D=0
M1348 258 468 466 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=80560 $D=0
M1349 259 469 467 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=85190 $D=0
M1350 468 81 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=80560 $D=0
M1351 469 81 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=85190 $D=0
M1352 8 82 470 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=80560 $D=0
M1353 8 82 471 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=85190 $D=0
M1354 472 83 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=80560 $D=0
M1355 473 83 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=85190 $D=0
M1356 474 470 244 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=80560 $D=0
M1357 475 471 245 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=85190 $D=0
M1358 8 474 765 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=80560 $D=0
M1359 8 475 766 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=85190 $D=0
M1360 476 765 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=80560 $D=0
M1361 477 766 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=85190 $D=0
M1362 474 82 476 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=80560 $D=0
M1363 475 82 477 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=85190 $D=0
M1364 476 472 254 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=80560 $D=0
M1365 477 473 255 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=85190 $D=0
M1366 258 478 476 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=80560 $D=0
M1367 259 479 477 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=85190 $D=0
M1368 478 84 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=80560 $D=0
M1369 479 84 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=85190 $D=0
M1370 8 85 480 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=80560 $D=0
M1371 8 85 481 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=85190 $D=0
M1372 482 86 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=80560 $D=0
M1373 483 86 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=85190 $D=0
M1374 484 480 244 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=80560 $D=0
M1375 485 481 245 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=85190 $D=0
M1376 8 484 767 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=80560 $D=0
M1377 8 485 768 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=85190 $D=0
M1378 486 767 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=80560 $D=0
M1379 487 768 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=85190 $D=0
M1380 484 85 486 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=80560 $D=0
M1381 485 85 487 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=85190 $D=0
M1382 486 482 254 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=80560 $D=0
M1383 487 483 255 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=85190 $D=0
M1384 258 488 486 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=80560 $D=0
M1385 259 489 487 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=85190 $D=0
M1386 488 87 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=80560 $D=0
M1387 489 87 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=85190 $D=0
M1388 8 88 490 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=80560 $D=0
M1389 8 88 491 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=85190 $D=0
M1390 492 89 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=80560 $D=0
M1391 493 89 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=85190 $D=0
M1392 494 490 244 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=80560 $D=0
M1393 495 491 245 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=85190 $D=0
M1394 8 494 769 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=80560 $D=0
M1395 8 495 770 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=85190 $D=0
M1396 496 769 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=80560 $D=0
M1397 497 770 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=85190 $D=0
M1398 494 88 496 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=80560 $D=0
M1399 495 88 497 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=85190 $D=0
M1400 496 492 254 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=80560 $D=0
M1401 497 493 255 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=85190 $D=0
M1402 258 498 496 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=80560 $D=0
M1403 259 499 497 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=85190 $D=0
M1404 498 90 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=80560 $D=0
M1405 499 90 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=85190 $D=0
M1406 8 91 500 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=80560 $D=0
M1407 8 91 501 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=85190 $D=0
M1408 502 92 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=80560 $D=0
M1409 503 92 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=85190 $D=0
M1410 504 500 244 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=80560 $D=0
M1411 505 501 245 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=85190 $D=0
M1412 8 504 771 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=80560 $D=0
M1413 8 505 772 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=85190 $D=0
M1414 506 771 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=80560 $D=0
M1415 507 772 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=85190 $D=0
M1416 504 91 506 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=80560 $D=0
M1417 505 91 507 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=85190 $D=0
M1418 506 502 254 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=80560 $D=0
M1419 507 503 255 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=85190 $D=0
M1420 258 508 506 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=80560 $D=0
M1421 259 509 507 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=85190 $D=0
M1422 508 93 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=80560 $D=0
M1423 509 93 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=85190 $D=0
M1424 8 94 510 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=80560 $D=0
M1425 8 94 511 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=85190 $D=0
M1426 512 95 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=80560 $D=0
M1427 513 95 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=85190 $D=0
M1428 514 510 244 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=80560 $D=0
M1429 515 511 245 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=85190 $D=0
M1430 8 514 773 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=80560 $D=0
M1431 8 515 774 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=85190 $D=0
M1432 516 773 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=80560 $D=0
M1433 517 774 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=85190 $D=0
M1434 514 94 516 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=80560 $D=0
M1435 515 94 517 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=85190 $D=0
M1436 516 512 254 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=80560 $D=0
M1437 517 513 255 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=85190 $D=0
M1438 258 518 516 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=80560 $D=0
M1439 259 519 517 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=85190 $D=0
M1440 518 96 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=80560 $D=0
M1441 519 96 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=85190 $D=0
M1442 8 97 520 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=80560 $D=0
M1443 8 97 521 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=85190 $D=0
M1444 522 98 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=80560 $D=0
M1445 523 98 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=85190 $D=0
M1446 524 520 244 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=80560 $D=0
M1447 525 521 245 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=85190 $D=0
M1448 8 524 775 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=80560 $D=0
M1449 8 525 776 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=85190 $D=0
M1450 526 775 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=80560 $D=0
M1451 527 776 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=85190 $D=0
M1452 524 97 526 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=80560 $D=0
M1453 525 97 527 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=85190 $D=0
M1454 526 522 254 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=80560 $D=0
M1455 527 523 255 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=85190 $D=0
M1456 258 528 526 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=80560 $D=0
M1457 259 529 527 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=85190 $D=0
M1458 528 99 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=80560 $D=0
M1459 529 99 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=85190 $D=0
M1460 8 100 530 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=80560 $D=0
M1461 8 100 531 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=85190 $D=0
M1462 532 101 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=80560 $D=0
M1463 533 101 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=85190 $D=0
M1464 534 530 244 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=80560 $D=0
M1465 535 531 245 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=85190 $D=0
M1466 8 534 777 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=80560 $D=0
M1467 8 535 778 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=85190 $D=0
M1468 536 777 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=80560 $D=0
M1469 537 778 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=85190 $D=0
M1470 534 100 536 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=80560 $D=0
M1471 535 100 537 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=85190 $D=0
M1472 536 532 254 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=80560 $D=0
M1473 537 533 255 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=85190 $D=0
M1474 258 538 536 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=80560 $D=0
M1475 259 539 537 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=85190 $D=0
M1476 538 102 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=80560 $D=0
M1477 539 102 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=85190 $D=0
M1478 8 103 540 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=80560 $D=0
M1479 8 103 541 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=85190 $D=0
M1480 542 104 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=80560 $D=0
M1481 543 104 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=85190 $D=0
M1482 544 540 244 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=80560 $D=0
M1483 545 541 245 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=85190 $D=0
M1484 8 544 779 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=80560 $D=0
M1485 8 545 780 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=85190 $D=0
M1486 546 779 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=80560 $D=0
M1487 547 780 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=85190 $D=0
M1488 544 103 546 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=80560 $D=0
M1489 545 103 547 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=85190 $D=0
M1490 546 542 254 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=80560 $D=0
M1491 547 543 255 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=85190 $D=0
M1492 258 548 546 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=80560 $D=0
M1493 259 549 547 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=85190 $D=0
M1494 548 105 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=80560 $D=0
M1495 549 105 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=85190 $D=0
M1496 8 106 550 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=80560 $D=0
M1497 8 106 551 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=85190 $D=0
M1498 552 107 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=80560 $D=0
M1499 553 107 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=85190 $D=0
M1500 554 550 244 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=80560 $D=0
M1501 555 551 245 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=85190 $D=0
M1502 8 554 781 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=80560 $D=0
M1503 8 555 782 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=85190 $D=0
M1504 556 781 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=80560 $D=0
M1505 557 782 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=85190 $D=0
M1506 554 106 556 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=80560 $D=0
M1507 555 106 557 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=85190 $D=0
M1508 556 552 254 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=80560 $D=0
M1509 557 553 255 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=85190 $D=0
M1510 258 558 556 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=80560 $D=0
M1511 259 559 557 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=85190 $D=0
M1512 558 108 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=80560 $D=0
M1513 559 108 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=85190 $D=0
M1514 8 109 560 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=80560 $D=0
M1515 8 109 561 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=85190 $D=0
M1516 562 110 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=80560 $D=0
M1517 563 110 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=85190 $D=0
M1518 5 562 254 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=80560 $D=0
M1519 5 563 255 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=85190 $D=0
M1520 258 560 5 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=80560 $D=0
M1521 259 561 5 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=85190 $D=0
M1522 8 566 564 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=80560 $D=0
M1523 8 567 565 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=85190 $D=0
M1524 566 111 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=80560 $D=0
M1525 567 111 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=85190 $D=0
M1526 783 254 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=80560 $D=0
M1527 784 255 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=85190 $D=0
M1528 568 566 783 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=80560 $D=0
M1529 569 567 784 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=85190 $D=0
M1530 8 568 570 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=80560 $D=0
M1531 8 569 571 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=85190 $D=0
M1532 785 570 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=80560 $D=0
M1533 786 571 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=85190 $D=0
M1534 568 564 785 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=80560 $D=0
M1535 569 565 786 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=85190 $D=0
M1536 8 575 573 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=80560 $D=0
M1537 8 576 574 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=85190 $D=0
M1538 575 111 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=80560 $D=0
M1539 576 111 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=85190 $D=0
M1540 787 258 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=80560 $D=0
M1541 788 259 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=85190 $D=0
M1542 577 575 787 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=80560 $D=0
M1543 578 576 788 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=85190 $D=0
M1544 8 577 117 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=80560 $D=0
M1545 8 578 118 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=85190 $D=0
M1546 789 117 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=80560 $D=0
M1547 790 118 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=85190 $D=0
M1548 577 573 789 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=80560 $D=0
M1549 578 574 790 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=85190 $D=0
M1550 579 119 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=80560 $D=0
M1551 580 119 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=85190 $D=0
M1552 581 119 570 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=80560 $D=0
M1553 582 119 571 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=85190 $D=0
M1554 121 579 581 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=80560 $D=0
M1555 122 580 582 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=85190 $D=0
M1556 583 123 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=80560 $D=0
M1557 584 123 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=85190 $D=0
M1558 585 123 117 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=80560 $D=0
M1559 586 123 118 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=85190 $D=0
M1560 791 583 585 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=80560 $D=0
M1561 792 584 586 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=85190 $D=0
M1562 8 117 791 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=80560 $D=0
M1563 8 118 792 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=85190 $D=0
M1564 587 125 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=80560 $D=0
M1565 588 125 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=85190 $D=0
M1566 589 125 585 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=80560 $D=0
M1567 590 125 586 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=85190 $D=0
M1568 10 587 589 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=80560 $D=0
M1569 11 588 590 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=85190 $D=0
M1570 592 591 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=80560 $D=0
M1571 593 126 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=85190 $D=0
M1572 8 596 594 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=80560 $D=0
M1573 8 597 595 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=85190 $D=0
M1574 598 581 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=80560 $D=0
M1575 599 582 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=85190 $D=0
M1576 596 581 591 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=80560 $D=0
M1577 597 582 126 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=85190 $D=0
M1578 592 598 596 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=80560 $D=0
M1579 593 599 597 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=85190 $D=0
M1580 600 594 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=80560 $D=0
M1581 601 595 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=85190 $D=0
M1582 128 594 589 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=80560 $D=0
M1583 591 595 590 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=85190 $D=0
M1584 581 600 128 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=80560 $D=0
M1585 582 601 591 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=85190 $D=0
M1586 602 128 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=80560 $D=0
M1587 603 591 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=85190 $D=0
M1588 604 594 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=80560 $D=0
M1589 605 595 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=85190 $D=0
M1590 606 594 602 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=80560 $D=0
M1591 607 595 603 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=85190 $D=0
M1592 589 604 606 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=80560 $D=0
M1593 590 605 607 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=85190 $D=0
M1594 803 581 8 8 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=80200 $D=0
M1595 804 582 8 8 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=84830 $D=0
M1596 608 589 803 8 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=80200 $D=0
M1597 609 590 804 8 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=84830 $D=0
M1598 610 606 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=80560 $D=0
M1599 611 607 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=85190 $D=0
M1600 612 581 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=80560 $D=0
M1601 613 582 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=85190 $D=0
M1602 8 589 612 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=80560 $D=0
M1603 8 590 613 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=85190 $D=0
M1604 614 581 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=80560 $D=0
M1605 615 582 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=85190 $D=0
M1606 8 589 614 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=80560 $D=0
M1607 8 590 615 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=85190 $D=0
M1608 805 581 8 8 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=80380 $D=0
M1609 806 582 8 8 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=85010 $D=0
M1610 618 589 805 8 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=80380 $D=0
M1611 619 590 806 8 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=85010 $D=0
M1612 8 614 618 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=80560 $D=0
M1613 8 615 619 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=85190 $D=0
M1614 620 129 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=80560 $D=0
M1615 621 129 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=85190 $D=0
M1616 622 129 608 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=80560 $D=0
M1617 623 129 609 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=85190 $D=0
M1618 612 620 622 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=80560 $D=0
M1619 613 621 623 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=85190 $D=0
M1620 624 129 610 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=80560 $D=0
M1621 625 129 611 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=85190 $D=0
M1622 618 620 624 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=80560 $D=0
M1623 619 621 625 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=85190 $D=0
M1624 626 130 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=80560 $D=0
M1625 627 130 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=85190 $D=0
M1626 628 130 624 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=80560 $D=0
M1627 629 130 625 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=85190 $D=0
M1628 622 626 628 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=80560 $D=0
M1629 623 627 629 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=85190 $D=0
M1630 12 628 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=80560 $D=0
M1631 13 629 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=85190 $D=0
M1632 630 131 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=80560 $D=0
M1633 631 131 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=85190 $D=0
M1634 632 131 132 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=80560 $D=0
M1635 633 131 133 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=85190 $D=0
M1636 134 630 632 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=80560 $D=0
M1637 135 631 633 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=85190 $D=0
M1638 634 131 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=80560 $D=0
M1639 635 131 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=85190 $D=0
M1640 636 131 136 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=80560 $D=0
M1641 637 131 137 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=85190 $D=0
M1642 138 634 636 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=80560 $D=0
M1643 139 635 637 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=85190 $D=0
M1644 638 131 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=80560 $D=0
M1645 639 131 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=85190 $D=0
M1646 640 131 140 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=80560 $D=0
M1647 641 131 141 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=85190 $D=0
M1648 113 638 640 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=80560 $D=0
M1649 115 639 641 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=85190 $D=0
M1650 642 131 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=80560 $D=0
M1651 643 131 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=85190 $D=0
M1652 644 131 142 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=80560 $D=0
M1653 645 131 143 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=85190 $D=0
M1654 114 642 644 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=80560 $D=0
M1655 116 643 645 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=85190 $D=0
M1656 646 131 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=80560 $D=0
M1657 647 131 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=85190 $D=0
M1658 648 131 5 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=80560 $D=0
M1659 649 131 5 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=85190 $D=0
M1660 144 646 648 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=80560 $D=0
M1661 145 647 649 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=85190 $D=0
M1662 8 581 793 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=80560 $D=0
M1663 8 582 794 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=85190 $D=0
M1664 135 793 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=80560 $D=0
M1665 132 794 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=85190 $D=0
M1666 650 146 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=80560 $D=0
M1667 651 146 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=85190 $D=0
M1668 147 146 135 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=80560 $D=0
M1669 148 146 132 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=85190 $D=0
M1670 632 650 147 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=80560 $D=0
M1671 633 651 148 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=85190 $D=0
M1672 652 149 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=80560 $D=0
M1673 653 149 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=85190 $D=0
M1674 120 149 147 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=80560 $D=0
M1675 124 149 148 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=85190 $D=0
M1676 636 652 120 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=80560 $D=0
M1677 637 653 124 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=85190 $D=0
M1678 654 150 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=80560 $D=0
M1679 655 150 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=85190 $D=0
M1680 112 150 120 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=80560 $D=0
M1681 127 150 124 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=85190 $D=0
M1682 640 654 112 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=80560 $D=0
M1683 641 655 127 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=85190 $D=0
M1684 656 151 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=80560 $D=0
M1685 657 151 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=85190 $D=0
M1686 152 151 112 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=80560 $D=0
M1687 153 151 127 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=85190 $D=0
M1688 644 656 152 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=80560 $D=0
M1689 645 657 153 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=85190 $D=0
M1690 658 154 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=80560 $D=0
M1691 659 154 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=85190 $D=0
M1692 230 154 152 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=80560 $D=0
M1693 231 154 153 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=85190 $D=0
M1694 648 658 230 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=80560 $D=0
M1695 649 659 231 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=85190 $D=0
M1696 660 155 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=80560 $D=0
M1697 661 155 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=85190 $D=0
M1698 662 155 117 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=80560 $D=0
M1699 663 155 118 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=85190 $D=0
M1700 10 660 662 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=80560 $D=0
M1701 11 661 663 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=85190 $D=0
M1702 664 570 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=80560 $D=0
M1703 665 571 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=85190 $D=0
M1704 8 662 664 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=80560 $D=0
M1705 8 663 665 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=85190 $D=0
M1706 807 570 8 8 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=80380 $D=0
M1707 808 571 8 8 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=85010 $D=0
M1708 668 662 807 8 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=80380 $D=0
M1709 669 663 808 8 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=85010 $D=0
M1710 8 664 668 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=80560 $D=0
M1711 8 665 669 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=85190 $D=0
M1712 795 156 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=80560 $D=0
M1713 796 670 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=85190 $D=0
M1714 8 668 795 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=80560 $D=0
M1715 8 669 796 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=85190 $D=0
M1716 670 795 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=80560 $D=0
M1717 157 796 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=85190 $D=0
M1718 809 570 8 8 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=80200 $D=0
M1719 810 571 8 8 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=84830 $D=0
M1720 671 673 809 8 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=80200 $D=0
M1721 672 674 810 8 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=84830 $D=0
M1722 673 662 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=80560 $D=0
M1723 674 663 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=85190 $D=0
M1724 675 671 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=80560 $D=0
M1725 676 672 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=85190 $D=0
M1726 8 156 675 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=80560 $D=0
M1727 8 670 676 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=85190 $D=0
M1728 678 158 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=80560 $D=0
M1729 679 677 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=85190 $D=0
M1730 677 675 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=80560 $D=0
M1731 159 676 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=85190 $D=0
M1732 8 678 677 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=80560 $D=0
M1733 8 679 159 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=85190 $D=0
M1734 681 680 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=80560 $D=0
M1735 682 160 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=85190 $D=0
M1736 8 685 683 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=80560 $D=0
M1737 8 686 684 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=85190 $D=0
M1738 687 121 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=80560 $D=0
M1739 688 122 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=85190 $D=0
M1740 685 121 680 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=80560 $D=0
M1741 686 122 160 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=85190 $D=0
M1742 681 687 685 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=80560 $D=0
M1743 682 688 686 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=85190 $D=0
M1744 689 683 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=80560 $D=0
M1745 690 684 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=85190 $D=0
M1746 161 683 5 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=80560 $D=0
M1747 680 684 5 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=85190 $D=0
M1748 121 689 161 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=80560 $D=0
M1749 122 690 680 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=85190 $D=0
M1750 691 161 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=80560 $D=0
M1751 692 680 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=85190 $D=0
M1752 693 683 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=80560 $D=0
M1753 694 684 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=85190 $D=0
M1754 232 683 691 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=80560 $D=0
M1755 233 684 692 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=85190 $D=0
M1756 5 693 232 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=80560 $D=0
M1757 5 694 233 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=85190 $D=0
M1758 695 162 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=80560 $D=0
M1759 696 162 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=85190 $D=0
M1760 697 162 232 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=80560 $D=0
M1761 698 162 233 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=85190 $D=0
M1762 12 695 697 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=80560 $D=0
M1763 13 696 698 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=85190 $D=0
M1764 699 163 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=80560 $D=0
M1765 700 163 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=85190 $D=0
M1766 701 163 697 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=80560 $D=0
M1767 702 163 698 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=85190 $D=0
M1768 5 699 701 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=80560 $D=0
M1769 5 700 702 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=85190 $D=0
M1770 703 111 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=80560 $D=0
M1771 704 111 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=85190 $D=0
M1772 8 703 705 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=80560 $D=0
M1773 8 704 706 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=85190 $D=0
M1774 707 111 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=80560 $D=0
M1775 708 111 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=85190 $D=0
M1776 709 705 701 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=80560 $D=0
M1777 710 706 702 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=85190 $D=0
M1778 8 709 797 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=80560 $D=0
M1779 8 710 798 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=85190 $D=0
M1780 711 797 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=80560 $D=0
M1781 712 798 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=85190 $D=0
M1782 709 703 711 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=80560 $D=0
M1783 710 704 712 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=85190 $D=0
M1784 713 707 711 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=80560 $D=0
M1785 714 708 712 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=85190 $D=0
M1786 8 717 715 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=80560 $D=0
M1787 8 718 716 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=85190 $D=0
M1788 717 111 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=80560 $D=0
M1789 718 111 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=85190 $D=0
M1790 799 713 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=80560 $D=0
M1791 800 714 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=85190 $D=0
M1792 719 717 799 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=80560 $D=0
M1793 720 718 800 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=85190 $D=0
M1794 8 719 121 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=80560 $D=0
M1795 8 720 122 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=85190 $D=0
M1796 801 121 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=80560 $D=0
M1797 802 122 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=85190 $D=0
M1798 719 715 801 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=80560 $D=0
M1799 720 716 802 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=85190 $D=0
.ENDS
***************************************
.SUBCKT ICV_31 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 129 130 131 132 133 134 135 136 137 138 139 140 141
+ 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161
+ 162 163 164 165
** N=824 EP=164 IP=1514 FDC=1800
M0 209 1 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=70050 $D=1
M1 210 1 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=74680 $D=1
M2 211 209 2 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=70050 $D=1
M3 212 210 3 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=74680 $D=1
M4 5 1 211 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=70050 $D=1
M5 5 1 212 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=74680 $D=1
M6 213 209 4 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=70050 $D=1
M7 214 210 4 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=74680 $D=1
M8 3 1 213 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=70050 $D=1
M9 3 1 214 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=74680 $D=1
M10 215 209 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=70050 $D=1
M11 216 210 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=74680 $D=1
M12 5 1 215 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=70050 $D=1
M13 3 1 216 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=74680 $D=1
M14 219 217 215 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=70050 $D=1
M15 220 218 216 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=74680 $D=1
M16 217 6 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=70050 $D=1
M17 218 6 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=74680 $D=1
M18 221 217 213 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=70050 $D=1
M19 222 218 214 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=74680 $D=1
M20 211 6 221 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=70050 $D=1
M21 212 6 222 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=74680 $D=1
M22 223 7 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=70050 $D=1
M23 224 7 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=74680 $D=1
M24 225 223 221 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=70050 $D=1
M25 226 224 222 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=74680 $D=1
M26 219 7 225 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=70050 $D=1
M27 220 7 226 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=74680 $D=1
M28 227 9 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=70050 $D=1
M29 228 9 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=74680 $D=1
M30 229 227 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=70050 $D=1
M31 230 228 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=74680 $D=1
M32 10 9 229 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=70050 $D=1
M33 11 9 230 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=74680 $D=1
M34 231 227 12 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=70050 $D=1
M35 232 228 13 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=74680 $D=1
M36 233 9 231 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=70050 $D=1
M37 234 9 232 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=74680 $D=1
M38 237 227 235 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=70050 $D=1
M39 238 228 236 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=74680 $D=1
M40 225 9 237 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=70050 $D=1
M41 226 9 238 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=74680 $D=1
M42 241 239 237 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=70050 $D=1
M43 242 240 238 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=74680 $D=1
M44 239 14 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=70050 $D=1
M45 240 14 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=74680 $D=1
M46 243 239 231 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=70050 $D=1
M47 244 240 232 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=74680 $D=1
M48 229 14 243 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=70050 $D=1
M49 230 14 244 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=74680 $D=1
M50 245 15 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=70050 $D=1
M51 246 15 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=74680 $D=1
M52 247 245 243 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=70050 $D=1
M53 248 246 244 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=74680 $D=1
M54 241 15 247 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=70050 $D=1
M55 242 15 248 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=74680 $D=1
M56 5 16 249 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=70050 $D=1
M57 5 16 250 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=74680 $D=1
M58 251 17 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=70050 $D=1
M59 252 17 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=74680 $D=1
M60 253 16 247 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=70050 $D=1
M61 254 16 248 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=74680 $D=1
M62 5 253 723 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=70050 $D=1
M63 5 254 724 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=74680 $D=1
M64 255 723 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=70050 $D=1
M65 256 724 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=74680 $D=1
M66 253 249 255 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=70050 $D=1
M67 254 250 256 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=74680 $D=1
M68 255 17 257 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=70050 $D=1
M69 256 17 258 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=74680 $D=1
M70 261 18 255 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=70050 $D=1
M71 262 18 256 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=74680 $D=1
M72 259 18 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=70050 $D=1
M73 260 18 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=74680 $D=1
M74 5 19 263 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=70050 $D=1
M75 5 19 264 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=74680 $D=1
M76 265 20 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=70050 $D=1
M77 266 20 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=74680 $D=1
M78 267 19 247 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=70050 $D=1
M79 268 19 248 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=74680 $D=1
M80 5 267 725 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=70050 $D=1
M81 5 268 726 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=74680 $D=1
M82 269 725 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=70050 $D=1
M83 270 726 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=74680 $D=1
M84 267 263 269 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=70050 $D=1
M85 268 264 270 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=74680 $D=1
M86 269 20 257 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=70050 $D=1
M87 270 20 258 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=74680 $D=1
M88 261 21 269 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=70050 $D=1
M89 262 21 270 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=74680 $D=1
M90 271 21 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=70050 $D=1
M91 272 21 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=74680 $D=1
M92 5 22 273 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=70050 $D=1
M93 5 22 274 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=74680 $D=1
M94 275 23 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=70050 $D=1
M95 276 23 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=74680 $D=1
M96 277 22 247 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=70050 $D=1
M97 278 22 248 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=74680 $D=1
M98 5 277 727 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=70050 $D=1
M99 5 278 728 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=74680 $D=1
M100 279 727 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=70050 $D=1
M101 280 728 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=74680 $D=1
M102 277 273 279 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=70050 $D=1
M103 278 274 280 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=74680 $D=1
M104 279 23 257 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=70050 $D=1
M105 280 23 258 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=74680 $D=1
M106 261 24 279 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=70050 $D=1
M107 262 24 280 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=74680 $D=1
M108 281 24 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=70050 $D=1
M109 282 24 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=74680 $D=1
M110 5 25 283 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=70050 $D=1
M111 5 25 284 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=74680 $D=1
M112 285 26 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=70050 $D=1
M113 286 26 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=74680 $D=1
M114 287 25 247 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=70050 $D=1
M115 288 25 248 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=74680 $D=1
M116 5 287 729 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=70050 $D=1
M117 5 288 730 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=74680 $D=1
M118 289 729 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=70050 $D=1
M119 290 730 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=74680 $D=1
M120 287 283 289 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=70050 $D=1
M121 288 284 290 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=74680 $D=1
M122 289 26 257 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=70050 $D=1
M123 290 26 258 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=74680 $D=1
M124 261 27 289 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=70050 $D=1
M125 262 27 290 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=74680 $D=1
M126 291 27 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=70050 $D=1
M127 292 27 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=74680 $D=1
M128 5 28 293 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=70050 $D=1
M129 5 28 294 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=74680 $D=1
M130 295 29 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=70050 $D=1
M131 296 29 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=74680 $D=1
M132 297 28 247 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=70050 $D=1
M133 298 28 248 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=74680 $D=1
M134 5 297 731 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=70050 $D=1
M135 5 298 732 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=74680 $D=1
M136 299 731 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=70050 $D=1
M137 300 732 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=74680 $D=1
M138 297 293 299 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=70050 $D=1
M139 298 294 300 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=74680 $D=1
M140 299 29 257 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=70050 $D=1
M141 300 29 258 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=74680 $D=1
M142 261 30 299 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=70050 $D=1
M143 262 30 300 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=74680 $D=1
M144 301 30 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=70050 $D=1
M145 302 30 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=74680 $D=1
M146 5 31 303 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=70050 $D=1
M147 5 31 304 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=74680 $D=1
M148 305 32 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=70050 $D=1
M149 306 32 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=74680 $D=1
M150 307 31 247 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=70050 $D=1
M151 308 31 248 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=74680 $D=1
M152 5 307 733 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=70050 $D=1
M153 5 308 734 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=74680 $D=1
M154 309 733 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=70050 $D=1
M155 310 734 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=74680 $D=1
M156 307 303 309 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=70050 $D=1
M157 308 304 310 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=74680 $D=1
M158 309 32 257 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=70050 $D=1
M159 310 32 258 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=74680 $D=1
M160 261 33 309 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=70050 $D=1
M161 262 33 310 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=74680 $D=1
M162 311 33 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=70050 $D=1
M163 312 33 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=74680 $D=1
M164 5 34 313 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=70050 $D=1
M165 5 34 314 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=74680 $D=1
M166 315 35 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=70050 $D=1
M167 316 35 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=74680 $D=1
M168 317 34 247 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=70050 $D=1
M169 318 34 248 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=74680 $D=1
M170 5 317 735 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=70050 $D=1
M171 5 318 736 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=74680 $D=1
M172 319 735 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=70050 $D=1
M173 320 736 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=74680 $D=1
M174 317 313 319 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=70050 $D=1
M175 318 314 320 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=74680 $D=1
M176 319 35 257 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=70050 $D=1
M177 320 35 258 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=74680 $D=1
M178 261 36 319 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=70050 $D=1
M179 262 36 320 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=74680 $D=1
M180 321 36 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=70050 $D=1
M181 322 36 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=74680 $D=1
M182 5 37 323 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=70050 $D=1
M183 5 37 324 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=74680 $D=1
M184 325 38 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=70050 $D=1
M185 326 38 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=74680 $D=1
M186 327 37 247 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=70050 $D=1
M187 328 37 248 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=74680 $D=1
M188 5 327 737 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=70050 $D=1
M189 5 328 738 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=74680 $D=1
M190 329 737 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=70050 $D=1
M191 330 738 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=74680 $D=1
M192 327 323 329 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=70050 $D=1
M193 328 324 330 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=74680 $D=1
M194 329 38 257 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=70050 $D=1
M195 330 38 258 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=74680 $D=1
M196 261 39 329 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=70050 $D=1
M197 262 39 330 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=74680 $D=1
M198 331 39 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=70050 $D=1
M199 332 39 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=74680 $D=1
M200 5 40 333 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=70050 $D=1
M201 5 40 334 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=74680 $D=1
M202 335 41 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=70050 $D=1
M203 336 41 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=74680 $D=1
M204 337 40 247 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=70050 $D=1
M205 338 40 248 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=74680 $D=1
M206 5 337 739 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=70050 $D=1
M207 5 338 740 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=74680 $D=1
M208 339 739 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=70050 $D=1
M209 340 740 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=74680 $D=1
M210 337 333 339 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=70050 $D=1
M211 338 334 340 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=74680 $D=1
M212 339 41 257 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=70050 $D=1
M213 340 41 258 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=74680 $D=1
M214 261 42 339 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=70050 $D=1
M215 262 42 340 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=74680 $D=1
M216 341 42 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=70050 $D=1
M217 342 42 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=74680 $D=1
M218 5 43 343 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=70050 $D=1
M219 5 43 344 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=74680 $D=1
M220 345 44 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=70050 $D=1
M221 346 44 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=74680 $D=1
M222 347 43 247 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=70050 $D=1
M223 348 43 248 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=74680 $D=1
M224 5 347 741 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=70050 $D=1
M225 5 348 742 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=74680 $D=1
M226 349 741 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=70050 $D=1
M227 350 742 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=74680 $D=1
M228 347 343 349 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=70050 $D=1
M229 348 344 350 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=74680 $D=1
M230 349 44 257 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=70050 $D=1
M231 350 44 258 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=74680 $D=1
M232 261 45 349 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=70050 $D=1
M233 262 45 350 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=74680 $D=1
M234 351 45 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=70050 $D=1
M235 352 45 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=74680 $D=1
M236 5 46 353 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=70050 $D=1
M237 5 46 354 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=74680 $D=1
M238 355 47 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=70050 $D=1
M239 356 47 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=74680 $D=1
M240 357 46 247 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=70050 $D=1
M241 358 46 248 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=74680 $D=1
M242 5 357 743 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=70050 $D=1
M243 5 358 744 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=74680 $D=1
M244 359 743 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=70050 $D=1
M245 360 744 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=74680 $D=1
M246 357 353 359 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=70050 $D=1
M247 358 354 360 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=74680 $D=1
M248 359 47 257 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=70050 $D=1
M249 360 47 258 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=74680 $D=1
M250 261 48 359 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=70050 $D=1
M251 262 48 360 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=74680 $D=1
M252 361 48 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=70050 $D=1
M253 362 48 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=74680 $D=1
M254 5 49 363 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=70050 $D=1
M255 5 49 364 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=74680 $D=1
M256 365 50 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=70050 $D=1
M257 366 50 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=74680 $D=1
M258 367 49 247 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=70050 $D=1
M259 368 49 248 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=74680 $D=1
M260 5 367 745 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=70050 $D=1
M261 5 368 746 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=74680 $D=1
M262 369 745 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=70050 $D=1
M263 370 746 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=74680 $D=1
M264 367 363 369 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=70050 $D=1
M265 368 364 370 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=74680 $D=1
M266 369 50 257 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=70050 $D=1
M267 370 50 258 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=74680 $D=1
M268 261 51 369 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=70050 $D=1
M269 262 51 370 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=74680 $D=1
M270 371 51 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=70050 $D=1
M271 372 51 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=74680 $D=1
M272 5 52 373 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=70050 $D=1
M273 5 52 374 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=74680 $D=1
M274 375 53 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=70050 $D=1
M275 376 53 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=74680 $D=1
M276 377 52 247 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=70050 $D=1
M277 378 52 248 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=74680 $D=1
M278 5 377 747 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=70050 $D=1
M279 5 378 748 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=74680 $D=1
M280 379 747 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=70050 $D=1
M281 380 748 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=74680 $D=1
M282 377 373 379 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=70050 $D=1
M283 378 374 380 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=74680 $D=1
M284 379 53 257 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=70050 $D=1
M285 380 53 258 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=74680 $D=1
M286 261 54 379 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=70050 $D=1
M287 262 54 380 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=74680 $D=1
M288 381 54 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=70050 $D=1
M289 382 54 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=74680 $D=1
M290 5 55 383 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=70050 $D=1
M291 5 55 384 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=74680 $D=1
M292 385 56 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=70050 $D=1
M293 386 56 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=74680 $D=1
M294 387 55 247 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=70050 $D=1
M295 388 55 248 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=74680 $D=1
M296 5 387 749 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=70050 $D=1
M297 5 388 750 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=74680 $D=1
M298 389 749 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=70050 $D=1
M299 390 750 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=74680 $D=1
M300 387 383 389 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=70050 $D=1
M301 388 384 390 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=74680 $D=1
M302 389 56 257 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=70050 $D=1
M303 390 56 258 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=74680 $D=1
M304 261 57 389 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=70050 $D=1
M305 262 57 390 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=74680 $D=1
M306 391 57 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=70050 $D=1
M307 392 57 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=74680 $D=1
M308 5 58 393 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=70050 $D=1
M309 5 58 394 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=74680 $D=1
M310 395 59 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=70050 $D=1
M311 396 59 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=74680 $D=1
M312 397 58 247 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=70050 $D=1
M313 398 58 248 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=74680 $D=1
M314 5 397 751 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=70050 $D=1
M315 5 398 752 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=74680 $D=1
M316 399 751 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=70050 $D=1
M317 400 752 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=74680 $D=1
M318 397 393 399 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=70050 $D=1
M319 398 394 400 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=74680 $D=1
M320 399 59 257 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=70050 $D=1
M321 400 59 258 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=74680 $D=1
M322 261 60 399 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=70050 $D=1
M323 262 60 400 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=74680 $D=1
M324 401 60 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=70050 $D=1
M325 402 60 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=74680 $D=1
M326 5 61 403 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=70050 $D=1
M327 5 61 404 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=74680 $D=1
M328 405 62 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=70050 $D=1
M329 406 62 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=74680 $D=1
M330 407 61 247 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=70050 $D=1
M331 408 61 248 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=74680 $D=1
M332 5 407 753 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=70050 $D=1
M333 5 408 754 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=74680 $D=1
M334 409 753 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=70050 $D=1
M335 410 754 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=74680 $D=1
M336 407 403 409 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=70050 $D=1
M337 408 404 410 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=74680 $D=1
M338 409 62 257 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=70050 $D=1
M339 410 62 258 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=74680 $D=1
M340 261 63 409 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=70050 $D=1
M341 262 63 410 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=74680 $D=1
M342 411 63 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=70050 $D=1
M343 412 63 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=74680 $D=1
M344 5 64 413 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=70050 $D=1
M345 5 64 414 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=74680 $D=1
M346 415 65 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=70050 $D=1
M347 416 65 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=74680 $D=1
M348 417 64 247 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=70050 $D=1
M349 418 64 248 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=74680 $D=1
M350 5 417 755 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=70050 $D=1
M351 5 418 756 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=74680 $D=1
M352 419 755 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=70050 $D=1
M353 420 756 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=74680 $D=1
M354 417 413 419 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=70050 $D=1
M355 418 414 420 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=74680 $D=1
M356 419 65 257 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=70050 $D=1
M357 420 65 258 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=74680 $D=1
M358 261 66 419 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=70050 $D=1
M359 262 66 420 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=74680 $D=1
M360 421 66 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=70050 $D=1
M361 422 66 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=74680 $D=1
M362 5 67 423 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=70050 $D=1
M363 5 67 424 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=74680 $D=1
M364 425 68 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=70050 $D=1
M365 426 68 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=74680 $D=1
M366 427 67 247 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=70050 $D=1
M367 428 67 248 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=74680 $D=1
M368 5 427 757 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=70050 $D=1
M369 5 428 758 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=74680 $D=1
M370 429 757 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=70050 $D=1
M371 430 758 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=74680 $D=1
M372 427 423 429 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=70050 $D=1
M373 428 424 430 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=74680 $D=1
M374 429 68 257 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=70050 $D=1
M375 430 68 258 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=74680 $D=1
M376 261 69 429 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=70050 $D=1
M377 262 69 430 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=74680 $D=1
M378 431 69 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=70050 $D=1
M379 432 69 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=74680 $D=1
M380 5 70 433 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=70050 $D=1
M381 5 70 434 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=74680 $D=1
M382 435 71 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=70050 $D=1
M383 436 71 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=74680 $D=1
M384 437 70 247 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=70050 $D=1
M385 438 70 248 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=74680 $D=1
M386 5 437 759 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=70050 $D=1
M387 5 438 760 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=74680 $D=1
M388 439 759 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=70050 $D=1
M389 440 760 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=74680 $D=1
M390 437 433 439 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=70050 $D=1
M391 438 434 440 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=74680 $D=1
M392 439 71 257 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=70050 $D=1
M393 440 71 258 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=74680 $D=1
M394 261 72 439 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=70050 $D=1
M395 262 72 440 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=74680 $D=1
M396 441 72 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=70050 $D=1
M397 442 72 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=74680 $D=1
M398 5 73 443 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=70050 $D=1
M399 5 73 444 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=74680 $D=1
M400 445 74 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=70050 $D=1
M401 446 74 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=74680 $D=1
M402 447 73 247 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=70050 $D=1
M403 448 73 248 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=74680 $D=1
M404 5 447 761 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=70050 $D=1
M405 5 448 762 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=74680 $D=1
M406 449 761 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=70050 $D=1
M407 450 762 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=74680 $D=1
M408 447 443 449 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=70050 $D=1
M409 448 444 450 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=74680 $D=1
M410 449 74 257 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=70050 $D=1
M411 450 74 258 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=74680 $D=1
M412 261 75 449 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=70050 $D=1
M413 262 75 450 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=74680 $D=1
M414 451 75 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=70050 $D=1
M415 452 75 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=74680 $D=1
M416 5 76 453 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=70050 $D=1
M417 5 76 454 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=74680 $D=1
M418 455 77 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=70050 $D=1
M419 456 77 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=74680 $D=1
M420 457 76 247 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=70050 $D=1
M421 458 76 248 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=74680 $D=1
M422 5 457 763 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=70050 $D=1
M423 5 458 764 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=74680 $D=1
M424 459 763 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=70050 $D=1
M425 460 764 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=74680 $D=1
M426 457 453 459 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=70050 $D=1
M427 458 454 460 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=74680 $D=1
M428 459 77 257 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=70050 $D=1
M429 460 77 258 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=74680 $D=1
M430 261 78 459 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=70050 $D=1
M431 262 78 460 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=74680 $D=1
M432 461 78 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=70050 $D=1
M433 462 78 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=74680 $D=1
M434 5 79 463 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=70050 $D=1
M435 5 79 464 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=74680 $D=1
M436 465 80 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=70050 $D=1
M437 466 80 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=74680 $D=1
M438 467 79 247 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=70050 $D=1
M439 468 79 248 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=74680 $D=1
M440 5 467 765 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=70050 $D=1
M441 5 468 766 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=74680 $D=1
M442 469 765 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=70050 $D=1
M443 470 766 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=74680 $D=1
M444 467 463 469 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=70050 $D=1
M445 468 464 470 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=74680 $D=1
M446 469 80 257 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=70050 $D=1
M447 470 80 258 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=74680 $D=1
M448 261 81 469 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=70050 $D=1
M449 262 81 470 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=74680 $D=1
M450 471 81 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=70050 $D=1
M451 472 81 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=74680 $D=1
M452 5 82 473 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=70050 $D=1
M453 5 82 474 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=74680 $D=1
M454 475 83 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=70050 $D=1
M455 476 83 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=74680 $D=1
M456 477 82 247 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=70050 $D=1
M457 478 82 248 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=74680 $D=1
M458 5 477 767 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=70050 $D=1
M459 5 478 768 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=74680 $D=1
M460 479 767 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=70050 $D=1
M461 480 768 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=74680 $D=1
M462 477 473 479 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=70050 $D=1
M463 478 474 480 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=74680 $D=1
M464 479 83 257 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=70050 $D=1
M465 480 83 258 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=74680 $D=1
M466 261 84 479 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=70050 $D=1
M467 262 84 480 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=74680 $D=1
M468 481 84 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=70050 $D=1
M469 482 84 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=74680 $D=1
M470 5 85 483 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=70050 $D=1
M471 5 85 484 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=74680 $D=1
M472 485 86 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=70050 $D=1
M473 486 86 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=74680 $D=1
M474 487 85 247 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=70050 $D=1
M475 488 85 248 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=74680 $D=1
M476 5 487 769 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=70050 $D=1
M477 5 488 770 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=74680 $D=1
M478 489 769 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=70050 $D=1
M479 490 770 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=74680 $D=1
M480 487 483 489 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=70050 $D=1
M481 488 484 490 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=74680 $D=1
M482 489 86 257 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=70050 $D=1
M483 490 86 258 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=74680 $D=1
M484 261 87 489 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=70050 $D=1
M485 262 87 490 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=74680 $D=1
M486 491 87 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=70050 $D=1
M487 492 87 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=74680 $D=1
M488 5 88 493 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=70050 $D=1
M489 5 88 494 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=74680 $D=1
M490 495 89 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=70050 $D=1
M491 496 89 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=74680 $D=1
M492 497 88 247 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=70050 $D=1
M493 498 88 248 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=74680 $D=1
M494 5 497 771 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=70050 $D=1
M495 5 498 772 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=74680 $D=1
M496 499 771 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=70050 $D=1
M497 500 772 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=74680 $D=1
M498 497 493 499 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=70050 $D=1
M499 498 494 500 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=74680 $D=1
M500 499 89 257 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=70050 $D=1
M501 500 89 258 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=74680 $D=1
M502 261 90 499 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=70050 $D=1
M503 262 90 500 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=74680 $D=1
M504 501 90 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=70050 $D=1
M505 502 90 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=74680 $D=1
M506 5 91 503 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=70050 $D=1
M507 5 91 504 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=74680 $D=1
M508 505 92 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=70050 $D=1
M509 506 92 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=74680 $D=1
M510 507 91 247 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=70050 $D=1
M511 508 91 248 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=74680 $D=1
M512 5 507 773 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=70050 $D=1
M513 5 508 774 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=74680 $D=1
M514 509 773 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=70050 $D=1
M515 510 774 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=74680 $D=1
M516 507 503 509 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=70050 $D=1
M517 508 504 510 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=74680 $D=1
M518 509 92 257 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=70050 $D=1
M519 510 92 258 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=74680 $D=1
M520 261 93 509 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=70050 $D=1
M521 262 93 510 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=74680 $D=1
M522 511 93 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=70050 $D=1
M523 512 93 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=74680 $D=1
M524 5 94 513 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=70050 $D=1
M525 5 94 514 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=74680 $D=1
M526 515 95 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=70050 $D=1
M527 516 95 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=74680 $D=1
M528 517 94 247 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=70050 $D=1
M529 518 94 248 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=74680 $D=1
M530 5 517 775 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=70050 $D=1
M531 5 518 776 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=74680 $D=1
M532 519 775 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=70050 $D=1
M533 520 776 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=74680 $D=1
M534 517 513 519 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=70050 $D=1
M535 518 514 520 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=74680 $D=1
M536 519 95 257 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=70050 $D=1
M537 520 95 258 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=74680 $D=1
M538 261 96 519 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=70050 $D=1
M539 262 96 520 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=74680 $D=1
M540 521 96 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=70050 $D=1
M541 522 96 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=74680 $D=1
M542 5 97 523 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=70050 $D=1
M543 5 97 524 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=74680 $D=1
M544 525 98 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=70050 $D=1
M545 526 98 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=74680 $D=1
M546 527 97 247 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=70050 $D=1
M547 528 97 248 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=74680 $D=1
M548 5 527 777 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=70050 $D=1
M549 5 528 778 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=74680 $D=1
M550 529 777 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=70050 $D=1
M551 530 778 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=74680 $D=1
M552 527 523 529 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=70050 $D=1
M553 528 524 530 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=74680 $D=1
M554 529 98 257 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=70050 $D=1
M555 530 98 258 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=74680 $D=1
M556 261 99 529 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=70050 $D=1
M557 262 99 530 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=74680 $D=1
M558 531 99 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=70050 $D=1
M559 532 99 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=74680 $D=1
M560 5 100 533 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=70050 $D=1
M561 5 100 534 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=74680 $D=1
M562 535 101 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=70050 $D=1
M563 536 101 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=74680 $D=1
M564 537 100 247 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=70050 $D=1
M565 538 100 248 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=74680 $D=1
M566 5 537 779 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=70050 $D=1
M567 5 538 780 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=74680 $D=1
M568 539 779 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=70050 $D=1
M569 540 780 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=74680 $D=1
M570 537 533 539 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=70050 $D=1
M571 538 534 540 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=74680 $D=1
M572 539 101 257 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=70050 $D=1
M573 540 101 258 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=74680 $D=1
M574 261 102 539 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=70050 $D=1
M575 262 102 540 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=74680 $D=1
M576 541 102 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=70050 $D=1
M577 542 102 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=74680 $D=1
M578 5 103 543 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=70050 $D=1
M579 5 103 544 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=74680 $D=1
M580 545 104 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=70050 $D=1
M581 546 104 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=74680 $D=1
M582 547 103 247 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=70050 $D=1
M583 548 103 248 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=74680 $D=1
M584 5 547 781 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=70050 $D=1
M585 5 548 782 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=74680 $D=1
M586 549 781 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=70050 $D=1
M587 550 782 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=74680 $D=1
M588 547 543 549 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=70050 $D=1
M589 548 544 550 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=74680 $D=1
M590 549 104 257 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=70050 $D=1
M591 550 104 258 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=74680 $D=1
M592 261 105 549 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=70050 $D=1
M593 262 105 550 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=74680 $D=1
M594 551 105 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=70050 $D=1
M595 552 105 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=74680 $D=1
M596 5 106 553 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=70050 $D=1
M597 5 106 554 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=74680 $D=1
M598 555 107 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=70050 $D=1
M599 556 107 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=74680 $D=1
M600 557 106 247 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=70050 $D=1
M601 558 106 248 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=74680 $D=1
M602 5 557 783 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=70050 $D=1
M603 5 558 784 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=74680 $D=1
M604 559 783 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=70050 $D=1
M605 560 784 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=74680 $D=1
M606 557 553 559 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=70050 $D=1
M607 558 554 560 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=74680 $D=1
M608 559 107 257 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=70050 $D=1
M609 560 107 258 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=74680 $D=1
M610 261 109 559 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=70050 $D=1
M611 262 109 560 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=74680 $D=1
M612 561 109 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=70050 $D=1
M613 562 109 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=74680 $D=1
M614 5 110 563 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=70050 $D=1
M615 5 110 564 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=74680 $D=1
M616 565 111 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=70050 $D=1
M617 566 111 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=74680 $D=1
M618 5 111 257 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=70050 $D=1
M619 5 111 258 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=74680 $D=1
M620 261 110 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=70050 $D=1
M621 262 110 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=74680 $D=1
M622 5 569 567 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=70050 $D=1
M623 5 570 568 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=74680 $D=1
M624 569 112 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=70050 $D=1
M625 570 112 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=74680 $D=1
M626 785 257 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=70050 $D=1
M627 786 258 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=74680 $D=1
M628 571 567 785 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=70050 $D=1
M629 572 568 786 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=74680 $D=1
M630 5 571 573 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=70050 $D=1
M631 5 572 574 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=74680 $D=1
M632 787 573 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=70050 $D=1
M633 788 574 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=74680 $D=1
M634 571 569 787 5 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=70050 $D=1
M635 572 570 788 5 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=74680 $D=1
M636 5 577 575 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=70050 $D=1
M637 5 578 576 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=74680 $D=1
M638 577 112 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=70050 $D=1
M639 578 112 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=74680 $D=1
M640 789 261 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=70050 $D=1
M641 790 262 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=74680 $D=1
M642 579 575 789 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=70050 $D=1
M643 580 576 790 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=74680 $D=1
M644 5 579 116 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=70050 $D=1
M645 5 580 117 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=74680 $D=1
M646 791 116 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=70050 $D=1
M647 792 117 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=74680 $D=1
M648 579 577 791 5 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=70050 $D=1
M649 580 578 792 5 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=74680 $D=1
M650 581 120 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=70050 $D=1
M651 582 120 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=74680 $D=1
M652 583 581 573 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=70050 $D=1
M653 584 582 574 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=74680 $D=1
M654 121 120 583 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=70050 $D=1
M655 122 120 584 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=74680 $D=1
M656 585 123 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=70050 $D=1
M657 586 123 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=74680 $D=1
M658 587 585 116 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=70050 $D=1
M659 588 586 117 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=74680 $D=1
M660 793 123 587 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=70050 $D=1
M661 794 123 588 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=74680 $D=1
M662 5 116 793 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=70050 $D=1
M663 5 117 794 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=74680 $D=1
M664 589 124 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=70050 $D=1
M665 590 124 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=74680 $D=1
M666 591 589 587 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=70050 $D=1
M667 592 590 588 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=74680 $D=1
M668 10 124 591 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=70050 $D=1
M669 11 124 592 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=74680 $D=1
M670 594 593 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=70050 $D=1
M671 595 125 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=74680 $D=1
M672 5 598 596 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=70050 $D=1
M673 5 599 597 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=74680 $D=1
M674 600 583 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=70050 $D=1
M675 601 584 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=74680 $D=1
M676 598 600 593 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=70050 $D=1
M677 599 601 125 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=74680 $D=1
M678 594 583 598 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=70050 $D=1
M679 595 584 599 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=74680 $D=1
M680 602 596 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=70050 $D=1
M681 603 597 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=74680 $D=1
M682 126 602 591 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=70050 $D=1
M683 593 603 592 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=74680 $D=1
M684 583 596 126 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=70050 $D=1
M685 584 597 593 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=74680 $D=1
M686 604 126 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=70050 $D=1
M687 605 593 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=74680 $D=1
M688 606 596 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=70050 $D=1
M689 607 597 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=74680 $D=1
M690 608 606 604 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=70050 $D=1
M691 609 607 605 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=74680 $D=1
M692 591 596 608 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=70050 $D=1
M693 592 597 609 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=74680 $D=1
M694 610 583 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=70050 $D=1
M695 611 584 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=74680 $D=1
M696 5 591 610 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=70050 $D=1
M697 5 592 611 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=74680 $D=1
M698 612 608 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=70050 $D=1
M699 613 609 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=74680 $D=1
M700 813 583 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=70050 $D=1
M701 814 584 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=74680 $D=1
M702 614 591 813 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=70050 $D=1
M703 615 592 814 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=74680 $D=1
M704 815 583 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=70050 $D=1
M705 816 584 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=74680 $D=1
M706 616 591 815 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=70050 $D=1
M707 617 592 816 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=74680 $D=1
M708 620 583 618 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=70050 $D=1
M709 621 584 619 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=74680 $D=1
M710 618 591 620 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=70050 $D=1
M711 619 592 621 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=74680 $D=1
M712 5 616 618 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=70050 $D=1
M713 5 617 619 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=74680 $D=1
M714 622 129 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=70050 $D=1
M715 623 129 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=74680 $D=1
M716 624 622 610 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=70050 $D=1
M717 625 623 611 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=74680 $D=1
M718 614 129 624 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=70050 $D=1
M719 615 129 625 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=74680 $D=1
M720 626 622 612 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=70050 $D=1
M721 627 623 613 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=74680 $D=1
M722 620 129 626 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=70050 $D=1
M723 621 129 627 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=74680 $D=1
M724 628 130 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=70050 $D=1
M725 629 130 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=74680 $D=1
M726 630 628 626 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=70050 $D=1
M727 631 629 627 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=74680 $D=1
M728 624 130 630 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=70050 $D=1
M729 625 130 631 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=74680 $D=1
M730 12 630 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=70050 $D=1
M731 13 631 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=74680 $D=1
M732 632 131 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=70050 $D=1
M733 633 131 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=74680 $D=1
M734 634 632 132 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=70050 $D=1
M735 635 633 133 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=74680 $D=1
M736 134 131 634 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=70050 $D=1
M737 135 131 635 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=74680 $D=1
M738 636 131 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=70050 $D=1
M739 637 131 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=74680 $D=1
M740 638 636 136 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=70050 $D=1
M741 639 637 137 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=74680 $D=1
M742 138 131 638 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=70050 $D=1
M743 139 131 639 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=74680 $D=1
M744 640 131 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=70050 $D=1
M745 641 131 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=74680 $D=1
M746 642 640 127 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=70050 $D=1
M747 643 641 140 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=74680 $D=1
M748 114 131 642 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=70050 $D=1
M749 115 131 643 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=74680 $D=1
M750 644 131 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=70050 $D=1
M751 645 131 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=74680 $D=1
M752 646 644 141 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=70050 $D=1
M753 647 645 142 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=74680 $D=1
M754 143 131 646 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=70050 $D=1
M755 144 131 647 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=74680 $D=1
M756 648 131 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=70050 $D=1
M757 649 131 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=74680 $D=1
M758 650 648 145 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=70050 $D=1
M759 651 649 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=74680 $D=1
M760 146 131 650 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=70050 $D=1
M761 147 131 651 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=74680 $D=1
M762 5 583 795 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=70050 $D=1
M763 5 584 796 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=74680 $D=1
M764 135 795 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=70050 $D=1
M765 132 796 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=74680 $D=1
M766 652 148 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=70050 $D=1
M767 653 148 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=74680 $D=1
M768 150 652 135 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=70050 $D=1
M769 151 653 132 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=74680 $D=1
M770 634 148 150 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=70050 $D=1
M771 635 148 151 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=74680 $D=1
M772 654 152 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=70050 $D=1
M773 655 152 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=74680 $D=1
M774 118 654 150 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=70050 $D=1
M775 119 655 151 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=74680 $D=1
M776 638 152 118 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=70050 $D=1
M777 639 152 119 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=74680 $D=1
M778 656 153 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=70050 $D=1
M779 657 153 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=74680 $D=1
M780 108 656 118 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=70050 $D=1
M781 113 657 119 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=74680 $D=1
M782 642 153 108 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=70050 $D=1
M783 643 153 113 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=74680 $D=1
M784 658 154 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=70050 $D=1
M785 659 154 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=74680 $D=1
M786 149 658 108 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=70050 $D=1
M787 155 659 113 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=74680 $D=1
M788 646 154 149 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=70050 $D=1
M789 647 154 155 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=74680 $D=1
M790 660 156 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=70050 $D=1
M791 661 156 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=74680 $D=1
M792 233 660 149 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=70050 $D=1
M793 234 661 155 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=74680 $D=1
M794 650 156 233 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=70050 $D=1
M795 651 156 234 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=74680 $D=1
M796 662 157 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=70050 $D=1
M797 663 157 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=74680 $D=1
M798 664 662 116 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=70050 $D=1
M799 665 663 117 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=74680 $D=1
M800 10 157 664 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=70050 $D=1
M801 11 157 665 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=74680 $D=1
M802 817 573 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=70050 $D=1
M803 818 574 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=74680 $D=1
M804 666 664 817 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=70050 $D=1
M805 667 665 818 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=74680 $D=1
M806 670 573 668 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=70050 $D=1
M807 671 574 669 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=74680 $D=1
M808 668 664 670 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=70050 $D=1
M809 669 665 671 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=74680 $D=1
M810 5 666 668 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=70050 $D=1
M811 5 667 669 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=74680 $D=1
M812 819 158 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=70050 $D=1
M813 820 672 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=74680 $D=1
M814 797 670 819 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=70050 $D=1
M815 798 671 820 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=74680 $D=1
M816 672 797 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=70050 $D=1
M817 159 798 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=74680 $D=1
M818 673 573 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=70050 $D=1
M819 674 574 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=74680 $D=1
M820 5 675 673 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=70050 $D=1
M821 5 676 674 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=74680 $D=1
M822 675 664 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=70050 $D=1
M823 676 665 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=74680 $D=1
M824 821 673 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=70050 $D=1
M825 822 674 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=74680 $D=1
M826 677 158 821 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=70050 $D=1
M827 678 672 822 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=74680 $D=1
M828 680 160 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=70050 $D=1
M829 681 679 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=74680 $D=1
M830 823 677 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=70050 $D=1
M831 824 678 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=74680 $D=1
M832 679 680 823 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=70050 $D=1
M833 161 681 824 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=74680 $D=1
M834 683 682 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=70050 $D=1
M835 684 162 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=74680 $D=1
M836 5 687 685 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=70050 $D=1
M837 5 688 686 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=74680 $D=1
M838 689 121 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=70050 $D=1
M839 690 122 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=74680 $D=1
M840 687 689 682 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=70050 $D=1
M841 688 690 162 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=74680 $D=1
M842 683 121 687 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=70050 $D=1
M843 684 122 688 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=74680 $D=1
M844 691 685 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=70050 $D=1
M845 692 686 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=74680 $D=1
M846 163 691 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=70050 $D=1
M847 682 692 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=74680 $D=1
M848 121 685 163 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=70050 $D=1
M849 122 686 682 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=74680 $D=1
M850 693 163 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=70050 $D=1
M851 694 682 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=74680 $D=1
M852 695 685 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=70050 $D=1
M853 696 686 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=74680 $D=1
M854 235 695 693 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=70050 $D=1
M855 236 696 694 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=74680 $D=1
M856 5 685 235 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=70050 $D=1
M857 5 686 236 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=74680 $D=1
M858 697 164 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=70050 $D=1
M859 698 164 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=74680 $D=1
M860 699 697 235 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=70050 $D=1
M861 700 698 236 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=74680 $D=1
M862 12 164 699 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=70050 $D=1
M863 13 164 700 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=74680 $D=1
M864 701 165 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=70050 $D=1
M865 702 165 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=74680 $D=1
M866 703 701 699 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=70050 $D=1
M867 704 702 700 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=74680 $D=1
M868 5 165 703 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=70050 $D=1
M869 5 165 704 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=74680 $D=1
M870 705 112 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=70050 $D=1
M871 706 112 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=74680 $D=1
M872 5 705 707 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=70050 $D=1
M873 5 706 708 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=74680 $D=1
M874 709 112 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=70050 $D=1
M875 710 112 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=74680 $D=1
M876 711 705 703 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=70050 $D=1
M877 712 706 704 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=74680 $D=1
M878 5 711 799 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=70050 $D=1
M879 5 712 800 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=74680 $D=1
M880 713 799 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=70050 $D=1
M881 714 800 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=74680 $D=1
M882 711 707 713 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=70050 $D=1
M883 712 708 714 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=74680 $D=1
M884 715 112 713 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=70050 $D=1
M885 716 112 714 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=74680 $D=1
M886 5 719 717 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=70050 $D=1
M887 5 720 718 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=74680 $D=1
M888 719 112 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=70050 $D=1
M889 720 112 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=74680 $D=1
M890 801 715 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=70050 $D=1
M891 802 716 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=74680 $D=1
M892 721 717 801 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=70050 $D=1
M893 722 718 802 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=74680 $D=1
M894 5 721 121 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=70050 $D=1
M895 5 722 122 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=74680 $D=1
M896 803 121 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=70050 $D=1
M897 804 122 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=74680 $D=1
M898 721 719 803 5 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=70050 $D=1
M899 722 720 804 5 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=74680 $D=1
M900 209 1 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=71300 $D=0
M901 210 1 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=75930 $D=0
M902 211 1 2 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=71300 $D=0
M903 212 1 3 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=75930 $D=0
M904 5 209 211 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=71300 $D=0
M905 5 210 212 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=75930 $D=0
M906 213 1 4 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=71300 $D=0
M907 214 1 4 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=75930 $D=0
M908 3 209 213 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=71300 $D=0
M909 3 210 214 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=75930 $D=0
M910 215 1 5 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=71300 $D=0
M911 216 1 5 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=75930 $D=0
M912 5 209 215 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=71300 $D=0
M913 3 210 216 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=75930 $D=0
M914 219 6 215 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=71300 $D=0
M915 220 6 216 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=75930 $D=0
M916 217 6 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=71300 $D=0
M917 218 6 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=75930 $D=0
M918 221 6 213 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=71300 $D=0
M919 222 6 214 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=75930 $D=0
M920 211 217 221 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=71300 $D=0
M921 212 218 222 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=75930 $D=0
M922 223 7 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=71300 $D=0
M923 224 7 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=75930 $D=0
M924 225 7 221 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=71300 $D=0
M925 226 7 222 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=75930 $D=0
M926 219 223 225 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=71300 $D=0
M927 220 224 226 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=75930 $D=0
M928 227 9 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=71300 $D=0
M929 228 9 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=75930 $D=0
M930 229 9 5 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=71300 $D=0
M931 230 9 5 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=75930 $D=0
M932 10 227 229 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=71300 $D=0
M933 11 228 230 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=75930 $D=0
M934 231 9 12 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=71300 $D=0
M935 232 9 13 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=75930 $D=0
M936 233 227 231 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=71300 $D=0
M937 234 228 232 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=75930 $D=0
M938 237 9 235 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=71300 $D=0
M939 238 9 236 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=75930 $D=0
M940 225 227 237 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=71300 $D=0
M941 226 228 238 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=75930 $D=0
M942 241 14 237 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=71300 $D=0
M943 242 14 238 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=75930 $D=0
M944 239 14 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=71300 $D=0
M945 240 14 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=75930 $D=0
M946 243 14 231 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=71300 $D=0
M947 244 14 232 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=75930 $D=0
M948 229 239 243 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=71300 $D=0
M949 230 240 244 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=75930 $D=0
M950 245 15 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=71300 $D=0
M951 246 15 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=75930 $D=0
M952 247 15 243 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=71300 $D=0
M953 248 15 244 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=75930 $D=0
M954 241 245 247 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=71300 $D=0
M955 242 246 248 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=75930 $D=0
M956 8 16 249 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=71300 $D=0
M957 8 16 250 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=75930 $D=0
M958 251 17 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=71300 $D=0
M959 252 17 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=75930 $D=0
M960 253 249 247 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=71300 $D=0
M961 254 250 248 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=75930 $D=0
M962 8 253 723 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=71300 $D=0
M963 8 254 724 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=75930 $D=0
M964 255 723 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=71300 $D=0
M965 256 724 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=75930 $D=0
M966 253 16 255 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=71300 $D=0
M967 254 16 256 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=75930 $D=0
M968 255 251 257 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=71300 $D=0
M969 256 252 258 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=75930 $D=0
M970 261 259 255 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=71300 $D=0
M971 262 260 256 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=75930 $D=0
M972 259 18 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=71300 $D=0
M973 260 18 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=75930 $D=0
M974 8 19 263 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=71300 $D=0
M975 8 19 264 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=75930 $D=0
M976 265 20 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=71300 $D=0
M977 266 20 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=75930 $D=0
M978 267 263 247 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=71300 $D=0
M979 268 264 248 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=75930 $D=0
M980 8 267 725 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=71300 $D=0
M981 8 268 726 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=75930 $D=0
M982 269 725 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=71300 $D=0
M983 270 726 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=75930 $D=0
M984 267 19 269 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=71300 $D=0
M985 268 19 270 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=75930 $D=0
M986 269 265 257 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=71300 $D=0
M987 270 266 258 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=75930 $D=0
M988 261 271 269 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=71300 $D=0
M989 262 272 270 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=75930 $D=0
M990 271 21 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=71300 $D=0
M991 272 21 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=75930 $D=0
M992 8 22 273 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=71300 $D=0
M993 8 22 274 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=75930 $D=0
M994 275 23 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=71300 $D=0
M995 276 23 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=75930 $D=0
M996 277 273 247 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=71300 $D=0
M997 278 274 248 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=75930 $D=0
M998 8 277 727 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=71300 $D=0
M999 8 278 728 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=75930 $D=0
M1000 279 727 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=71300 $D=0
M1001 280 728 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=75930 $D=0
M1002 277 22 279 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=71300 $D=0
M1003 278 22 280 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=75930 $D=0
M1004 279 275 257 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=71300 $D=0
M1005 280 276 258 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=75930 $D=0
M1006 261 281 279 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=71300 $D=0
M1007 262 282 280 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=75930 $D=0
M1008 281 24 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=71300 $D=0
M1009 282 24 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=75930 $D=0
M1010 8 25 283 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=71300 $D=0
M1011 8 25 284 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=75930 $D=0
M1012 285 26 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=71300 $D=0
M1013 286 26 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=75930 $D=0
M1014 287 283 247 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=71300 $D=0
M1015 288 284 248 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=75930 $D=0
M1016 8 287 729 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=71300 $D=0
M1017 8 288 730 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=75930 $D=0
M1018 289 729 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=71300 $D=0
M1019 290 730 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=75930 $D=0
M1020 287 25 289 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=71300 $D=0
M1021 288 25 290 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=75930 $D=0
M1022 289 285 257 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=71300 $D=0
M1023 290 286 258 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=75930 $D=0
M1024 261 291 289 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=71300 $D=0
M1025 262 292 290 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=75930 $D=0
M1026 291 27 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=71300 $D=0
M1027 292 27 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=75930 $D=0
M1028 8 28 293 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=71300 $D=0
M1029 8 28 294 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=75930 $D=0
M1030 295 29 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=71300 $D=0
M1031 296 29 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=75930 $D=0
M1032 297 293 247 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=71300 $D=0
M1033 298 294 248 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=75930 $D=0
M1034 8 297 731 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=71300 $D=0
M1035 8 298 732 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=75930 $D=0
M1036 299 731 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=71300 $D=0
M1037 300 732 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=75930 $D=0
M1038 297 28 299 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=71300 $D=0
M1039 298 28 300 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=75930 $D=0
M1040 299 295 257 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=71300 $D=0
M1041 300 296 258 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=75930 $D=0
M1042 261 301 299 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=71300 $D=0
M1043 262 302 300 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=75930 $D=0
M1044 301 30 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=71300 $D=0
M1045 302 30 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=75930 $D=0
M1046 8 31 303 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=71300 $D=0
M1047 8 31 304 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=75930 $D=0
M1048 305 32 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=71300 $D=0
M1049 306 32 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=75930 $D=0
M1050 307 303 247 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=71300 $D=0
M1051 308 304 248 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=75930 $D=0
M1052 8 307 733 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=71300 $D=0
M1053 8 308 734 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=75930 $D=0
M1054 309 733 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=71300 $D=0
M1055 310 734 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=75930 $D=0
M1056 307 31 309 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=71300 $D=0
M1057 308 31 310 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=75930 $D=0
M1058 309 305 257 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=71300 $D=0
M1059 310 306 258 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=75930 $D=0
M1060 261 311 309 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=71300 $D=0
M1061 262 312 310 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=75930 $D=0
M1062 311 33 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=71300 $D=0
M1063 312 33 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=75930 $D=0
M1064 8 34 313 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=71300 $D=0
M1065 8 34 314 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=75930 $D=0
M1066 315 35 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=71300 $D=0
M1067 316 35 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=75930 $D=0
M1068 317 313 247 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=71300 $D=0
M1069 318 314 248 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=75930 $D=0
M1070 8 317 735 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=71300 $D=0
M1071 8 318 736 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=75930 $D=0
M1072 319 735 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=71300 $D=0
M1073 320 736 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=75930 $D=0
M1074 317 34 319 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=71300 $D=0
M1075 318 34 320 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=75930 $D=0
M1076 319 315 257 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=71300 $D=0
M1077 320 316 258 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=75930 $D=0
M1078 261 321 319 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=71300 $D=0
M1079 262 322 320 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=75930 $D=0
M1080 321 36 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=71300 $D=0
M1081 322 36 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=75930 $D=0
M1082 8 37 323 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=71300 $D=0
M1083 8 37 324 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=75930 $D=0
M1084 325 38 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=71300 $D=0
M1085 326 38 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=75930 $D=0
M1086 327 323 247 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=71300 $D=0
M1087 328 324 248 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=75930 $D=0
M1088 8 327 737 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=71300 $D=0
M1089 8 328 738 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=75930 $D=0
M1090 329 737 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=71300 $D=0
M1091 330 738 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=75930 $D=0
M1092 327 37 329 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=71300 $D=0
M1093 328 37 330 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=75930 $D=0
M1094 329 325 257 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=71300 $D=0
M1095 330 326 258 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=75930 $D=0
M1096 261 331 329 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=71300 $D=0
M1097 262 332 330 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=75930 $D=0
M1098 331 39 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=71300 $D=0
M1099 332 39 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=75930 $D=0
M1100 8 40 333 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=71300 $D=0
M1101 8 40 334 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=75930 $D=0
M1102 335 41 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=71300 $D=0
M1103 336 41 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=75930 $D=0
M1104 337 333 247 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=71300 $D=0
M1105 338 334 248 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=75930 $D=0
M1106 8 337 739 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=71300 $D=0
M1107 8 338 740 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=75930 $D=0
M1108 339 739 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=71300 $D=0
M1109 340 740 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=75930 $D=0
M1110 337 40 339 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=71300 $D=0
M1111 338 40 340 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=75930 $D=0
M1112 339 335 257 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=71300 $D=0
M1113 340 336 258 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=75930 $D=0
M1114 261 341 339 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=71300 $D=0
M1115 262 342 340 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=75930 $D=0
M1116 341 42 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=71300 $D=0
M1117 342 42 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=75930 $D=0
M1118 8 43 343 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=71300 $D=0
M1119 8 43 344 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=75930 $D=0
M1120 345 44 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=71300 $D=0
M1121 346 44 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=75930 $D=0
M1122 347 343 247 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=71300 $D=0
M1123 348 344 248 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=75930 $D=0
M1124 8 347 741 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=71300 $D=0
M1125 8 348 742 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=75930 $D=0
M1126 349 741 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=71300 $D=0
M1127 350 742 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=75930 $D=0
M1128 347 43 349 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=71300 $D=0
M1129 348 43 350 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=75930 $D=0
M1130 349 345 257 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=71300 $D=0
M1131 350 346 258 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=75930 $D=0
M1132 261 351 349 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=71300 $D=0
M1133 262 352 350 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=75930 $D=0
M1134 351 45 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=71300 $D=0
M1135 352 45 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=75930 $D=0
M1136 8 46 353 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=71300 $D=0
M1137 8 46 354 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=75930 $D=0
M1138 355 47 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=71300 $D=0
M1139 356 47 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=75930 $D=0
M1140 357 353 247 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=71300 $D=0
M1141 358 354 248 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=75930 $D=0
M1142 8 357 743 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=71300 $D=0
M1143 8 358 744 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=75930 $D=0
M1144 359 743 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=71300 $D=0
M1145 360 744 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=75930 $D=0
M1146 357 46 359 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=71300 $D=0
M1147 358 46 360 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=75930 $D=0
M1148 359 355 257 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=71300 $D=0
M1149 360 356 258 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=75930 $D=0
M1150 261 361 359 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=71300 $D=0
M1151 262 362 360 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=75930 $D=0
M1152 361 48 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=71300 $D=0
M1153 362 48 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=75930 $D=0
M1154 8 49 363 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=71300 $D=0
M1155 8 49 364 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=75930 $D=0
M1156 365 50 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=71300 $D=0
M1157 366 50 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=75930 $D=0
M1158 367 363 247 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=71300 $D=0
M1159 368 364 248 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=75930 $D=0
M1160 8 367 745 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=71300 $D=0
M1161 8 368 746 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=75930 $D=0
M1162 369 745 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=71300 $D=0
M1163 370 746 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=75930 $D=0
M1164 367 49 369 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=71300 $D=0
M1165 368 49 370 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=75930 $D=0
M1166 369 365 257 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=71300 $D=0
M1167 370 366 258 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=75930 $D=0
M1168 261 371 369 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=71300 $D=0
M1169 262 372 370 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=75930 $D=0
M1170 371 51 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=71300 $D=0
M1171 372 51 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=75930 $D=0
M1172 8 52 373 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=71300 $D=0
M1173 8 52 374 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=75930 $D=0
M1174 375 53 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=71300 $D=0
M1175 376 53 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=75930 $D=0
M1176 377 373 247 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=71300 $D=0
M1177 378 374 248 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=75930 $D=0
M1178 8 377 747 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=71300 $D=0
M1179 8 378 748 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=75930 $D=0
M1180 379 747 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=71300 $D=0
M1181 380 748 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=75930 $D=0
M1182 377 52 379 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=71300 $D=0
M1183 378 52 380 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=75930 $D=0
M1184 379 375 257 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=71300 $D=0
M1185 380 376 258 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=75930 $D=0
M1186 261 381 379 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=71300 $D=0
M1187 262 382 380 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=75930 $D=0
M1188 381 54 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=71300 $D=0
M1189 382 54 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=75930 $D=0
M1190 8 55 383 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=71300 $D=0
M1191 8 55 384 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=75930 $D=0
M1192 385 56 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=71300 $D=0
M1193 386 56 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=75930 $D=0
M1194 387 383 247 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=71300 $D=0
M1195 388 384 248 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=75930 $D=0
M1196 8 387 749 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=71300 $D=0
M1197 8 388 750 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=75930 $D=0
M1198 389 749 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=71300 $D=0
M1199 390 750 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=75930 $D=0
M1200 387 55 389 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=71300 $D=0
M1201 388 55 390 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=75930 $D=0
M1202 389 385 257 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=71300 $D=0
M1203 390 386 258 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=75930 $D=0
M1204 261 391 389 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=71300 $D=0
M1205 262 392 390 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=75930 $D=0
M1206 391 57 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=71300 $D=0
M1207 392 57 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=75930 $D=0
M1208 8 58 393 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=71300 $D=0
M1209 8 58 394 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=75930 $D=0
M1210 395 59 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=71300 $D=0
M1211 396 59 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=75930 $D=0
M1212 397 393 247 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=71300 $D=0
M1213 398 394 248 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=75930 $D=0
M1214 8 397 751 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=71300 $D=0
M1215 8 398 752 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=75930 $D=0
M1216 399 751 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=71300 $D=0
M1217 400 752 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=75930 $D=0
M1218 397 58 399 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=71300 $D=0
M1219 398 58 400 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=75930 $D=0
M1220 399 395 257 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=71300 $D=0
M1221 400 396 258 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=75930 $D=0
M1222 261 401 399 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=71300 $D=0
M1223 262 402 400 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=75930 $D=0
M1224 401 60 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=71300 $D=0
M1225 402 60 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=75930 $D=0
M1226 8 61 403 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=71300 $D=0
M1227 8 61 404 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=75930 $D=0
M1228 405 62 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=71300 $D=0
M1229 406 62 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=75930 $D=0
M1230 407 403 247 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=71300 $D=0
M1231 408 404 248 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=75930 $D=0
M1232 8 407 753 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=71300 $D=0
M1233 8 408 754 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=75930 $D=0
M1234 409 753 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=71300 $D=0
M1235 410 754 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=75930 $D=0
M1236 407 61 409 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=71300 $D=0
M1237 408 61 410 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=75930 $D=0
M1238 409 405 257 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=71300 $D=0
M1239 410 406 258 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=75930 $D=0
M1240 261 411 409 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=71300 $D=0
M1241 262 412 410 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=75930 $D=0
M1242 411 63 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=71300 $D=0
M1243 412 63 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=75930 $D=0
M1244 8 64 413 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=71300 $D=0
M1245 8 64 414 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=75930 $D=0
M1246 415 65 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=71300 $D=0
M1247 416 65 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=75930 $D=0
M1248 417 413 247 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=71300 $D=0
M1249 418 414 248 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=75930 $D=0
M1250 8 417 755 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=71300 $D=0
M1251 8 418 756 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=75930 $D=0
M1252 419 755 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=71300 $D=0
M1253 420 756 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=75930 $D=0
M1254 417 64 419 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=71300 $D=0
M1255 418 64 420 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=75930 $D=0
M1256 419 415 257 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=71300 $D=0
M1257 420 416 258 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=75930 $D=0
M1258 261 421 419 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=71300 $D=0
M1259 262 422 420 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=75930 $D=0
M1260 421 66 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=71300 $D=0
M1261 422 66 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=75930 $D=0
M1262 8 67 423 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=71300 $D=0
M1263 8 67 424 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=75930 $D=0
M1264 425 68 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=71300 $D=0
M1265 426 68 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=75930 $D=0
M1266 427 423 247 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=71300 $D=0
M1267 428 424 248 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=75930 $D=0
M1268 8 427 757 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=71300 $D=0
M1269 8 428 758 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=75930 $D=0
M1270 429 757 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=71300 $D=0
M1271 430 758 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=75930 $D=0
M1272 427 67 429 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=71300 $D=0
M1273 428 67 430 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=75930 $D=0
M1274 429 425 257 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=71300 $D=0
M1275 430 426 258 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=75930 $D=0
M1276 261 431 429 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=71300 $D=0
M1277 262 432 430 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=75930 $D=0
M1278 431 69 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=71300 $D=0
M1279 432 69 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=75930 $D=0
M1280 8 70 433 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=71300 $D=0
M1281 8 70 434 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=75930 $D=0
M1282 435 71 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=71300 $D=0
M1283 436 71 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=75930 $D=0
M1284 437 433 247 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=71300 $D=0
M1285 438 434 248 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=75930 $D=0
M1286 8 437 759 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=71300 $D=0
M1287 8 438 760 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=75930 $D=0
M1288 439 759 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=71300 $D=0
M1289 440 760 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=75930 $D=0
M1290 437 70 439 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=71300 $D=0
M1291 438 70 440 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=75930 $D=0
M1292 439 435 257 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=71300 $D=0
M1293 440 436 258 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=75930 $D=0
M1294 261 441 439 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=71300 $D=0
M1295 262 442 440 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=75930 $D=0
M1296 441 72 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=71300 $D=0
M1297 442 72 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=75930 $D=0
M1298 8 73 443 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=71300 $D=0
M1299 8 73 444 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=75930 $D=0
M1300 445 74 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=71300 $D=0
M1301 446 74 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=75930 $D=0
M1302 447 443 247 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=71300 $D=0
M1303 448 444 248 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=75930 $D=0
M1304 8 447 761 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=71300 $D=0
M1305 8 448 762 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=75930 $D=0
M1306 449 761 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=71300 $D=0
M1307 450 762 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=75930 $D=0
M1308 447 73 449 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=71300 $D=0
M1309 448 73 450 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=75930 $D=0
M1310 449 445 257 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=71300 $D=0
M1311 450 446 258 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=75930 $D=0
M1312 261 451 449 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=71300 $D=0
M1313 262 452 450 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=75930 $D=0
M1314 451 75 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=71300 $D=0
M1315 452 75 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=75930 $D=0
M1316 8 76 453 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=71300 $D=0
M1317 8 76 454 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=75930 $D=0
M1318 455 77 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=71300 $D=0
M1319 456 77 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=75930 $D=0
M1320 457 453 247 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=71300 $D=0
M1321 458 454 248 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=75930 $D=0
M1322 8 457 763 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=71300 $D=0
M1323 8 458 764 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=75930 $D=0
M1324 459 763 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=71300 $D=0
M1325 460 764 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=75930 $D=0
M1326 457 76 459 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=71300 $D=0
M1327 458 76 460 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=75930 $D=0
M1328 459 455 257 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=71300 $D=0
M1329 460 456 258 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=75930 $D=0
M1330 261 461 459 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=71300 $D=0
M1331 262 462 460 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=75930 $D=0
M1332 461 78 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=71300 $D=0
M1333 462 78 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=75930 $D=0
M1334 8 79 463 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=71300 $D=0
M1335 8 79 464 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=75930 $D=0
M1336 465 80 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=71300 $D=0
M1337 466 80 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=75930 $D=0
M1338 467 463 247 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=71300 $D=0
M1339 468 464 248 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=75930 $D=0
M1340 8 467 765 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=71300 $D=0
M1341 8 468 766 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=75930 $D=0
M1342 469 765 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=71300 $D=0
M1343 470 766 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=75930 $D=0
M1344 467 79 469 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=71300 $D=0
M1345 468 79 470 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=75930 $D=0
M1346 469 465 257 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=71300 $D=0
M1347 470 466 258 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=75930 $D=0
M1348 261 471 469 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=71300 $D=0
M1349 262 472 470 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=75930 $D=0
M1350 471 81 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=71300 $D=0
M1351 472 81 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=75930 $D=0
M1352 8 82 473 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=71300 $D=0
M1353 8 82 474 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=75930 $D=0
M1354 475 83 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=71300 $D=0
M1355 476 83 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=75930 $D=0
M1356 477 473 247 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=71300 $D=0
M1357 478 474 248 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=75930 $D=0
M1358 8 477 767 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=71300 $D=0
M1359 8 478 768 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=75930 $D=0
M1360 479 767 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=71300 $D=0
M1361 480 768 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=75930 $D=0
M1362 477 82 479 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=71300 $D=0
M1363 478 82 480 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=75930 $D=0
M1364 479 475 257 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=71300 $D=0
M1365 480 476 258 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=75930 $D=0
M1366 261 481 479 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=71300 $D=0
M1367 262 482 480 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=75930 $D=0
M1368 481 84 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=71300 $D=0
M1369 482 84 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=75930 $D=0
M1370 8 85 483 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=71300 $D=0
M1371 8 85 484 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=75930 $D=0
M1372 485 86 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=71300 $D=0
M1373 486 86 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=75930 $D=0
M1374 487 483 247 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=71300 $D=0
M1375 488 484 248 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=75930 $D=0
M1376 8 487 769 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=71300 $D=0
M1377 8 488 770 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=75930 $D=0
M1378 489 769 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=71300 $D=0
M1379 490 770 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=75930 $D=0
M1380 487 85 489 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=71300 $D=0
M1381 488 85 490 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=75930 $D=0
M1382 489 485 257 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=71300 $D=0
M1383 490 486 258 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=75930 $D=0
M1384 261 491 489 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=71300 $D=0
M1385 262 492 490 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=75930 $D=0
M1386 491 87 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=71300 $D=0
M1387 492 87 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=75930 $D=0
M1388 8 88 493 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=71300 $D=0
M1389 8 88 494 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=75930 $D=0
M1390 495 89 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=71300 $D=0
M1391 496 89 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=75930 $D=0
M1392 497 493 247 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=71300 $D=0
M1393 498 494 248 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=75930 $D=0
M1394 8 497 771 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=71300 $D=0
M1395 8 498 772 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=75930 $D=0
M1396 499 771 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=71300 $D=0
M1397 500 772 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=75930 $D=0
M1398 497 88 499 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=71300 $D=0
M1399 498 88 500 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=75930 $D=0
M1400 499 495 257 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=71300 $D=0
M1401 500 496 258 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=75930 $D=0
M1402 261 501 499 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=71300 $D=0
M1403 262 502 500 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=75930 $D=0
M1404 501 90 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=71300 $D=0
M1405 502 90 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=75930 $D=0
M1406 8 91 503 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=71300 $D=0
M1407 8 91 504 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=75930 $D=0
M1408 505 92 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=71300 $D=0
M1409 506 92 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=75930 $D=0
M1410 507 503 247 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=71300 $D=0
M1411 508 504 248 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=75930 $D=0
M1412 8 507 773 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=71300 $D=0
M1413 8 508 774 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=75930 $D=0
M1414 509 773 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=71300 $D=0
M1415 510 774 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=75930 $D=0
M1416 507 91 509 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=71300 $D=0
M1417 508 91 510 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=75930 $D=0
M1418 509 505 257 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=71300 $D=0
M1419 510 506 258 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=75930 $D=0
M1420 261 511 509 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=71300 $D=0
M1421 262 512 510 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=75930 $D=0
M1422 511 93 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=71300 $D=0
M1423 512 93 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=75930 $D=0
M1424 8 94 513 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=71300 $D=0
M1425 8 94 514 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=75930 $D=0
M1426 515 95 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=71300 $D=0
M1427 516 95 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=75930 $D=0
M1428 517 513 247 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=71300 $D=0
M1429 518 514 248 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=75930 $D=0
M1430 8 517 775 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=71300 $D=0
M1431 8 518 776 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=75930 $D=0
M1432 519 775 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=71300 $D=0
M1433 520 776 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=75930 $D=0
M1434 517 94 519 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=71300 $D=0
M1435 518 94 520 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=75930 $D=0
M1436 519 515 257 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=71300 $D=0
M1437 520 516 258 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=75930 $D=0
M1438 261 521 519 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=71300 $D=0
M1439 262 522 520 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=75930 $D=0
M1440 521 96 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=71300 $D=0
M1441 522 96 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=75930 $D=0
M1442 8 97 523 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=71300 $D=0
M1443 8 97 524 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=75930 $D=0
M1444 525 98 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=71300 $D=0
M1445 526 98 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=75930 $D=0
M1446 527 523 247 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=71300 $D=0
M1447 528 524 248 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=75930 $D=0
M1448 8 527 777 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=71300 $D=0
M1449 8 528 778 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=75930 $D=0
M1450 529 777 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=71300 $D=0
M1451 530 778 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=75930 $D=0
M1452 527 97 529 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=71300 $D=0
M1453 528 97 530 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=75930 $D=0
M1454 529 525 257 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=71300 $D=0
M1455 530 526 258 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=75930 $D=0
M1456 261 531 529 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=71300 $D=0
M1457 262 532 530 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=75930 $D=0
M1458 531 99 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=71300 $D=0
M1459 532 99 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=75930 $D=0
M1460 8 100 533 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=71300 $D=0
M1461 8 100 534 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=75930 $D=0
M1462 535 101 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=71300 $D=0
M1463 536 101 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=75930 $D=0
M1464 537 533 247 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=71300 $D=0
M1465 538 534 248 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=75930 $D=0
M1466 8 537 779 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=71300 $D=0
M1467 8 538 780 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=75930 $D=0
M1468 539 779 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=71300 $D=0
M1469 540 780 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=75930 $D=0
M1470 537 100 539 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=71300 $D=0
M1471 538 100 540 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=75930 $D=0
M1472 539 535 257 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=71300 $D=0
M1473 540 536 258 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=75930 $D=0
M1474 261 541 539 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=71300 $D=0
M1475 262 542 540 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=75930 $D=0
M1476 541 102 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=71300 $D=0
M1477 542 102 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=75930 $D=0
M1478 8 103 543 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=71300 $D=0
M1479 8 103 544 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=75930 $D=0
M1480 545 104 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=71300 $D=0
M1481 546 104 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=75930 $D=0
M1482 547 543 247 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=71300 $D=0
M1483 548 544 248 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=75930 $D=0
M1484 8 547 781 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=71300 $D=0
M1485 8 548 782 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=75930 $D=0
M1486 549 781 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=71300 $D=0
M1487 550 782 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=75930 $D=0
M1488 547 103 549 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=71300 $D=0
M1489 548 103 550 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=75930 $D=0
M1490 549 545 257 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=71300 $D=0
M1491 550 546 258 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=75930 $D=0
M1492 261 551 549 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=71300 $D=0
M1493 262 552 550 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=75930 $D=0
M1494 551 105 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=71300 $D=0
M1495 552 105 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=75930 $D=0
M1496 8 106 553 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=71300 $D=0
M1497 8 106 554 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=75930 $D=0
M1498 555 107 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=71300 $D=0
M1499 556 107 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=75930 $D=0
M1500 557 553 247 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=71300 $D=0
M1501 558 554 248 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=75930 $D=0
M1502 8 557 783 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=71300 $D=0
M1503 8 558 784 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=75930 $D=0
M1504 559 783 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=71300 $D=0
M1505 560 784 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=75930 $D=0
M1506 557 106 559 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=71300 $D=0
M1507 558 106 560 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=75930 $D=0
M1508 559 555 257 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=71300 $D=0
M1509 560 556 258 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=75930 $D=0
M1510 261 561 559 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=71300 $D=0
M1511 262 562 560 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=75930 $D=0
M1512 561 109 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=71300 $D=0
M1513 562 109 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=75930 $D=0
M1514 8 110 563 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=71300 $D=0
M1515 8 110 564 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=75930 $D=0
M1516 565 111 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=71300 $D=0
M1517 566 111 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=75930 $D=0
M1518 5 565 257 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=71300 $D=0
M1519 5 566 258 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=75930 $D=0
M1520 261 563 5 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=71300 $D=0
M1521 262 564 5 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=75930 $D=0
M1522 8 569 567 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=71300 $D=0
M1523 8 570 568 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=75930 $D=0
M1524 569 112 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=71300 $D=0
M1525 570 112 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=75930 $D=0
M1526 785 257 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=71300 $D=0
M1527 786 258 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=75930 $D=0
M1528 571 569 785 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=71300 $D=0
M1529 572 570 786 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=75930 $D=0
M1530 8 571 573 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=71300 $D=0
M1531 8 572 574 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=75930 $D=0
M1532 787 573 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=71300 $D=0
M1533 788 574 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=75930 $D=0
M1534 571 567 787 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=71300 $D=0
M1535 572 568 788 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=75930 $D=0
M1536 8 577 575 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=71300 $D=0
M1537 8 578 576 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=75930 $D=0
M1538 577 112 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=71300 $D=0
M1539 578 112 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=75930 $D=0
M1540 789 261 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=71300 $D=0
M1541 790 262 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=75930 $D=0
M1542 579 577 789 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=71300 $D=0
M1543 580 578 790 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=75930 $D=0
M1544 8 579 116 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=71300 $D=0
M1545 8 580 117 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=75930 $D=0
M1546 791 116 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=71300 $D=0
M1547 792 117 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=75930 $D=0
M1548 579 575 791 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=71300 $D=0
M1549 580 576 792 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=75930 $D=0
M1550 581 120 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=71300 $D=0
M1551 582 120 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=75930 $D=0
M1552 583 120 573 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=71300 $D=0
M1553 584 120 574 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=75930 $D=0
M1554 121 581 583 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=71300 $D=0
M1555 122 582 584 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=75930 $D=0
M1556 585 123 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=71300 $D=0
M1557 586 123 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=75930 $D=0
M1558 587 123 116 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=71300 $D=0
M1559 588 123 117 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=75930 $D=0
M1560 793 585 587 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=71300 $D=0
M1561 794 586 588 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=75930 $D=0
M1562 8 116 793 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=71300 $D=0
M1563 8 117 794 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=75930 $D=0
M1564 589 124 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=71300 $D=0
M1565 590 124 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=75930 $D=0
M1566 591 124 587 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=71300 $D=0
M1567 592 124 588 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=75930 $D=0
M1568 10 589 591 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=71300 $D=0
M1569 11 590 592 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=75930 $D=0
M1570 594 593 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=71300 $D=0
M1571 595 125 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=75930 $D=0
M1572 8 598 596 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=71300 $D=0
M1573 8 599 597 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=75930 $D=0
M1574 600 583 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=71300 $D=0
M1575 601 584 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=75930 $D=0
M1576 598 583 593 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=71300 $D=0
M1577 599 584 125 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=75930 $D=0
M1578 594 600 598 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=71300 $D=0
M1579 595 601 599 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=75930 $D=0
M1580 602 596 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=71300 $D=0
M1581 603 597 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=75930 $D=0
M1582 126 596 591 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=71300 $D=0
M1583 593 597 592 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=75930 $D=0
M1584 583 602 126 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=71300 $D=0
M1585 584 603 593 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=75930 $D=0
M1586 604 126 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=71300 $D=0
M1587 605 593 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=75930 $D=0
M1588 606 596 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=71300 $D=0
M1589 607 597 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=75930 $D=0
M1590 608 596 604 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=71300 $D=0
M1591 609 597 605 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=75930 $D=0
M1592 591 606 608 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=71300 $D=0
M1593 592 607 609 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=75930 $D=0
M1594 805 583 8 8 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=70940 $D=0
M1595 806 584 8 8 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=75570 $D=0
M1596 610 591 805 8 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=70940 $D=0
M1597 611 592 806 8 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=75570 $D=0
M1598 612 608 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=71300 $D=0
M1599 613 609 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=75930 $D=0
M1600 614 583 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=71300 $D=0
M1601 615 584 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=75930 $D=0
M1602 8 591 614 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=71300 $D=0
M1603 8 592 615 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=75930 $D=0
M1604 616 583 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=71300 $D=0
M1605 617 584 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=75930 $D=0
M1606 8 591 616 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=71300 $D=0
M1607 8 592 617 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=75930 $D=0
M1608 807 583 8 8 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=71120 $D=0
M1609 808 584 8 8 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=75750 $D=0
M1610 620 591 807 8 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=71120 $D=0
M1611 621 592 808 8 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=75750 $D=0
M1612 8 616 620 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=71300 $D=0
M1613 8 617 621 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=75930 $D=0
M1614 622 129 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=71300 $D=0
M1615 623 129 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=75930 $D=0
M1616 624 129 610 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=71300 $D=0
M1617 625 129 611 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=75930 $D=0
M1618 614 622 624 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=71300 $D=0
M1619 615 623 625 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=75930 $D=0
M1620 626 129 612 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=71300 $D=0
M1621 627 129 613 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=75930 $D=0
M1622 620 622 626 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=71300 $D=0
M1623 621 623 627 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=75930 $D=0
M1624 628 130 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=71300 $D=0
M1625 629 130 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=75930 $D=0
M1626 630 130 626 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=71300 $D=0
M1627 631 130 627 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=75930 $D=0
M1628 624 628 630 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=71300 $D=0
M1629 625 629 631 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=75930 $D=0
M1630 12 630 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=71300 $D=0
M1631 13 631 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=75930 $D=0
M1632 632 131 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=71300 $D=0
M1633 633 131 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=75930 $D=0
M1634 634 131 132 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=71300 $D=0
M1635 635 131 133 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=75930 $D=0
M1636 134 632 634 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=71300 $D=0
M1637 135 633 635 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=75930 $D=0
M1638 636 131 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=71300 $D=0
M1639 637 131 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=75930 $D=0
M1640 638 131 136 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=71300 $D=0
M1641 639 131 137 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=75930 $D=0
M1642 138 636 638 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=71300 $D=0
M1643 139 637 639 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=75930 $D=0
M1644 640 131 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=71300 $D=0
M1645 641 131 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=75930 $D=0
M1646 642 131 127 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=71300 $D=0
M1647 643 131 140 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=75930 $D=0
M1648 114 640 642 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=71300 $D=0
M1649 115 641 643 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=75930 $D=0
M1650 644 131 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=71300 $D=0
M1651 645 131 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=75930 $D=0
M1652 646 131 141 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=71300 $D=0
M1653 647 131 142 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=75930 $D=0
M1654 143 644 646 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=71300 $D=0
M1655 144 645 647 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=75930 $D=0
M1656 648 131 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=71300 $D=0
M1657 649 131 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=75930 $D=0
M1658 650 131 145 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=71300 $D=0
M1659 651 131 5 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=75930 $D=0
M1660 146 648 650 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=71300 $D=0
M1661 147 649 651 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=75930 $D=0
M1662 8 583 795 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=71300 $D=0
M1663 8 584 796 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=75930 $D=0
M1664 135 795 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=71300 $D=0
M1665 132 796 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=75930 $D=0
M1666 652 148 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=71300 $D=0
M1667 653 148 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=75930 $D=0
M1668 150 148 135 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=71300 $D=0
M1669 151 148 132 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=75930 $D=0
M1670 634 652 150 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=71300 $D=0
M1671 635 653 151 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=75930 $D=0
M1672 654 152 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=71300 $D=0
M1673 655 152 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=75930 $D=0
M1674 118 152 150 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=71300 $D=0
M1675 119 152 151 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=75930 $D=0
M1676 638 654 118 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=71300 $D=0
M1677 639 655 119 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=75930 $D=0
M1678 656 153 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=71300 $D=0
M1679 657 153 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=75930 $D=0
M1680 108 153 118 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=71300 $D=0
M1681 113 153 119 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=75930 $D=0
M1682 642 656 108 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=71300 $D=0
M1683 643 657 113 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=75930 $D=0
M1684 658 154 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=71300 $D=0
M1685 659 154 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=75930 $D=0
M1686 149 154 108 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=71300 $D=0
M1687 155 154 113 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=75930 $D=0
M1688 646 658 149 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=71300 $D=0
M1689 647 659 155 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=75930 $D=0
M1690 660 156 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=71300 $D=0
M1691 661 156 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=75930 $D=0
M1692 233 156 149 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=71300 $D=0
M1693 234 156 155 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=75930 $D=0
M1694 650 660 233 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=71300 $D=0
M1695 651 661 234 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=75930 $D=0
M1696 662 157 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=71300 $D=0
M1697 663 157 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=75930 $D=0
M1698 664 157 116 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=71300 $D=0
M1699 665 157 117 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=75930 $D=0
M1700 10 662 664 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=71300 $D=0
M1701 11 663 665 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=75930 $D=0
M1702 666 573 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=71300 $D=0
M1703 667 574 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=75930 $D=0
M1704 8 664 666 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=71300 $D=0
M1705 8 665 667 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=75930 $D=0
M1706 809 573 8 8 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=71120 $D=0
M1707 810 574 8 8 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=75750 $D=0
M1708 670 664 809 8 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=71120 $D=0
M1709 671 665 810 8 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=75750 $D=0
M1710 8 666 670 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=71300 $D=0
M1711 8 667 671 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=75930 $D=0
M1712 797 158 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=71300 $D=0
M1713 798 672 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=75930 $D=0
M1714 8 670 797 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=71300 $D=0
M1715 8 671 798 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=75930 $D=0
M1716 672 797 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=71300 $D=0
M1717 159 798 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=75930 $D=0
M1718 811 573 8 8 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=70940 $D=0
M1719 812 574 8 8 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=75570 $D=0
M1720 673 675 811 8 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=70940 $D=0
M1721 674 676 812 8 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=75570 $D=0
M1722 675 664 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=71300 $D=0
M1723 676 665 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=75930 $D=0
M1724 677 673 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=71300 $D=0
M1725 678 674 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=75930 $D=0
M1726 8 158 677 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=71300 $D=0
M1727 8 672 678 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=75930 $D=0
M1728 680 160 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=71300 $D=0
M1729 681 679 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=75930 $D=0
M1730 679 677 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=71300 $D=0
M1731 161 678 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=75930 $D=0
M1732 8 680 679 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=71300 $D=0
M1733 8 681 161 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=75930 $D=0
M1734 683 682 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=71300 $D=0
M1735 684 162 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=75930 $D=0
M1736 8 687 685 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=71300 $D=0
M1737 8 688 686 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=75930 $D=0
M1738 689 121 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=71300 $D=0
M1739 690 122 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=75930 $D=0
M1740 687 121 682 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=71300 $D=0
M1741 688 122 162 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=75930 $D=0
M1742 683 689 687 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=71300 $D=0
M1743 684 690 688 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=75930 $D=0
M1744 691 685 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=71300 $D=0
M1745 692 686 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=75930 $D=0
M1746 163 685 5 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=71300 $D=0
M1747 682 686 5 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=75930 $D=0
M1748 121 691 163 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=71300 $D=0
M1749 122 692 682 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=75930 $D=0
M1750 693 163 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=71300 $D=0
M1751 694 682 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=75930 $D=0
M1752 695 685 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=71300 $D=0
M1753 696 686 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=75930 $D=0
M1754 235 685 693 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=71300 $D=0
M1755 236 686 694 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=75930 $D=0
M1756 5 695 235 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=71300 $D=0
M1757 5 696 236 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=75930 $D=0
M1758 697 164 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=71300 $D=0
M1759 698 164 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=75930 $D=0
M1760 699 164 235 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=71300 $D=0
M1761 700 164 236 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=75930 $D=0
M1762 12 697 699 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=71300 $D=0
M1763 13 698 700 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=75930 $D=0
M1764 701 165 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=71300 $D=0
M1765 702 165 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=75930 $D=0
M1766 703 165 699 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=71300 $D=0
M1767 704 165 700 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=75930 $D=0
M1768 5 701 703 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=71300 $D=0
M1769 5 702 704 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=75930 $D=0
M1770 705 112 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=71300 $D=0
M1771 706 112 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=75930 $D=0
M1772 8 705 707 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=71300 $D=0
M1773 8 706 708 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=75930 $D=0
M1774 709 112 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=71300 $D=0
M1775 710 112 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=75930 $D=0
M1776 711 707 703 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=71300 $D=0
M1777 712 708 704 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=75930 $D=0
M1778 8 711 799 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=71300 $D=0
M1779 8 712 800 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=75930 $D=0
M1780 713 799 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=71300 $D=0
M1781 714 800 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=75930 $D=0
M1782 711 705 713 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=71300 $D=0
M1783 712 706 714 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=75930 $D=0
M1784 715 709 713 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=71300 $D=0
M1785 716 710 714 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=75930 $D=0
M1786 8 719 717 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=71300 $D=0
M1787 8 720 718 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=75930 $D=0
M1788 719 112 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=71300 $D=0
M1789 720 112 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=75930 $D=0
M1790 801 715 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=71300 $D=0
M1791 802 716 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=75930 $D=0
M1792 721 719 801 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=71300 $D=0
M1793 722 720 802 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=75930 $D=0
M1794 8 721 121 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=71300 $D=0
M1795 8 722 122 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=75930 $D=0
M1796 803 121 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=71300 $D=0
M1797 804 122 8 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=75930 $D=0
M1798 721 717 803 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=71300 $D=0
M1799 722 718 804 8 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=75930 $D=0
.ENDS
***************************************
.SUBCKT ICV_32
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_33
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_34
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_35
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_36 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180
+ 181 182 183 184 185 186 187 188 189 190 191 192 193
** N=1461 EP=193 IP=2964 FDC=3600
M0 224 1 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=51530 $D=1
M1 225 1 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=56160 $D=1
M2 226 1 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=60790 $D=1
M3 227 1 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=65420 $D=1
M4 228 224 2 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=51530 $D=1
M5 229 225 3 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=56160 $D=1
M6 230 226 4 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=60790 $D=1
M7 231 227 5 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=65420 $D=1
M8 8 1 228 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=51530 $D=1
M9 8 1 229 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=56160 $D=1
M10 8 1 230 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=60790 $D=1
M11 8 1 231 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=65420 $D=1
M12 232 224 6 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=51530 $D=1
M13 233 225 6 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=56160 $D=1
M14 234 226 6 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=60790 $D=1
M15 235 227 6 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=65420 $D=1
M16 7 1 232 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=51530 $D=1
M17 7 1 233 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=56160 $D=1
M18 7 1 234 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=60790 $D=1
M19 7 1 235 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=65420 $D=1
M20 236 224 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=51530 $D=1
M21 237 225 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=56160 $D=1
M22 238 226 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=60790 $D=1
M23 239 227 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=65420 $D=1
M24 8 1 236 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=51530 $D=1
M25 8 1 237 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=56160 $D=1
M26 8 1 238 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=60790 $D=1
M27 8 1 239 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=65420 $D=1
M28 244 240 236 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=51530 $D=1
M29 245 241 237 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=56160 $D=1
M30 246 242 238 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=60790 $D=1
M31 247 243 239 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=65420 $D=1
M32 240 9 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=51530 $D=1
M33 241 9 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=56160 $D=1
M34 242 9 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=60790 $D=1
M35 243 9 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=65420 $D=1
M36 248 240 232 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=51530 $D=1
M37 249 241 233 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=56160 $D=1
M38 250 242 234 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=60790 $D=1
M39 251 243 235 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=65420 $D=1
M40 228 9 248 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=51530 $D=1
M41 229 9 249 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=56160 $D=1
M42 230 9 250 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=60790 $D=1
M43 231 9 251 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=65420 $D=1
M44 252 10 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=51530 $D=1
M45 253 10 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=56160 $D=1
M46 254 10 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=60790 $D=1
M47 255 10 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=65420 $D=1
M48 256 252 248 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=51530 $D=1
M49 257 253 249 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=56160 $D=1
M50 258 254 250 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=60790 $D=1
M51 259 255 251 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=65420 $D=1
M52 244 10 256 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=51530 $D=1
M53 245 10 257 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=56160 $D=1
M54 246 10 258 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=60790 $D=1
M55 247 10 259 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=65420 $D=1
M56 260 12 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=51530 $D=1
M57 261 12 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=56160 $D=1
M58 262 12 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=60790 $D=1
M59 263 12 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=65420 $D=1
M60 264 260 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=51530 $D=1
M61 265 261 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=56160 $D=1
M62 266 262 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=60790 $D=1
M63 267 263 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=65420 $D=1
M64 13 12 264 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=51530 $D=1
M65 14 12 265 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=56160 $D=1
M66 15 12 266 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=60790 $D=1
M67 16 12 267 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=65420 $D=1
M68 268 260 17 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=51530 $D=1
M69 269 261 18 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=56160 $D=1
M70 270 262 19 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=60790 $D=1
M71 271 263 20 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=65420 $D=1
M72 272 12 268 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=51530 $D=1
M73 273 12 269 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=56160 $D=1
M74 274 12 270 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=60790 $D=1
M75 275 12 271 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=65420 $D=1
M76 280 260 276 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=51530 $D=1
M77 281 261 277 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=56160 $D=1
M78 282 262 278 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=60790 $D=1
M79 283 263 279 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=65420 $D=1
M80 256 12 280 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=51530 $D=1
M81 257 12 281 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=56160 $D=1
M82 258 12 282 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=60790 $D=1
M83 259 12 283 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=65420 $D=1
M84 288 284 280 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=51530 $D=1
M85 289 285 281 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=56160 $D=1
M86 290 286 282 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=60790 $D=1
M87 291 287 283 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=65420 $D=1
M88 284 21 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=51530 $D=1
M89 285 21 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=56160 $D=1
M90 286 21 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=60790 $D=1
M91 287 21 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=65420 $D=1
M92 292 284 268 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=51530 $D=1
M93 293 285 269 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=56160 $D=1
M94 294 286 270 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=60790 $D=1
M95 295 287 271 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=65420 $D=1
M96 264 21 292 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=51530 $D=1
M97 265 21 293 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=56160 $D=1
M98 266 21 294 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=60790 $D=1
M99 267 21 295 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=65420 $D=1
M100 296 22 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=51530 $D=1
M101 297 22 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=56160 $D=1
M102 298 22 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=60790 $D=1
M103 299 22 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=65420 $D=1
M104 300 296 292 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=51530 $D=1
M105 301 297 293 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=56160 $D=1
M106 302 298 294 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=60790 $D=1
M107 303 299 295 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=65420 $D=1
M108 288 22 300 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=51530 $D=1
M109 289 22 301 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=56160 $D=1
M110 290 22 302 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=60790 $D=1
M111 291 22 303 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=65420 $D=1
M112 8 23 304 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=51530 $D=1
M113 8 23 305 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=56160 $D=1
M114 8 23 306 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=60790 $D=1
M115 8 23 307 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=65420 $D=1
M116 308 24 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=51530 $D=1
M117 309 24 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=56160 $D=1
M118 310 24 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=60790 $D=1
M119 311 24 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=65420 $D=1
M120 312 23 300 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=51530 $D=1
M121 313 23 301 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=56160 $D=1
M122 314 23 302 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=60790 $D=1
M123 315 23 303 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=65420 $D=1
M124 8 312 1258 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=51530 $D=1
M125 8 313 1259 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=56160 $D=1
M126 8 314 1260 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=60790 $D=1
M127 8 315 1261 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=65420 $D=1
M128 316 1258 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=51530 $D=1
M129 317 1259 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=56160 $D=1
M130 318 1260 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=60790 $D=1
M131 319 1261 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=65420 $D=1
M132 312 304 316 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=51530 $D=1
M133 313 305 317 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=56160 $D=1
M134 314 306 318 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=60790 $D=1
M135 315 307 319 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=65420 $D=1
M136 316 24 320 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=51530 $D=1
M137 317 24 321 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=56160 $D=1
M138 318 24 322 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=60790 $D=1
M139 319 24 323 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=65420 $D=1
M140 328 25 316 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=51530 $D=1
M141 329 25 317 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=56160 $D=1
M142 330 25 318 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=60790 $D=1
M143 331 25 319 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=65420 $D=1
M144 324 25 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=51530 $D=1
M145 325 25 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=56160 $D=1
M146 326 25 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=60790 $D=1
M147 327 25 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=65420 $D=1
M148 8 26 332 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=51530 $D=1
M149 8 26 333 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=56160 $D=1
M150 8 26 334 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=60790 $D=1
M151 8 26 335 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=65420 $D=1
M152 336 27 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=51530 $D=1
M153 337 27 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=56160 $D=1
M154 338 27 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=60790 $D=1
M155 339 27 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=65420 $D=1
M156 340 26 300 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=51530 $D=1
M157 341 26 301 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=56160 $D=1
M158 342 26 302 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=60790 $D=1
M159 343 26 303 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=65420 $D=1
M160 8 340 1262 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=51530 $D=1
M161 8 341 1263 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=56160 $D=1
M162 8 342 1264 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=60790 $D=1
M163 8 343 1265 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=65420 $D=1
M164 344 1262 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=51530 $D=1
M165 345 1263 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=56160 $D=1
M166 346 1264 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=60790 $D=1
M167 347 1265 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=65420 $D=1
M168 340 332 344 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=51530 $D=1
M169 341 333 345 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=56160 $D=1
M170 342 334 346 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=60790 $D=1
M171 343 335 347 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=65420 $D=1
M172 344 27 320 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=51530 $D=1
M173 345 27 321 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=56160 $D=1
M174 346 27 322 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=60790 $D=1
M175 347 27 323 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=65420 $D=1
M176 328 28 344 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=51530 $D=1
M177 329 28 345 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=56160 $D=1
M178 330 28 346 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=60790 $D=1
M179 331 28 347 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=65420 $D=1
M180 348 28 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=51530 $D=1
M181 349 28 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=56160 $D=1
M182 350 28 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=60790 $D=1
M183 351 28 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=65420 $D=1
M184 8 29 352 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=51530 $D=1
M185 8 29 353 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=56160 $D=1
M186 8 29 354 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=60790 $D=1
M187 8 29 355 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=65420 $D=1
M188 356 30 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=51530 $D=1
M189 357 30 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=56160 $D=1
M190 358 30 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=60790 $D=1
M191 359 30 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=65420 $D=1
M192 360 29 300 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=51530 $D=1
M193 361 29 301 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=56160 $D=1
M194 362 29 302 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=60790 $D=1
M195 363 29 303 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=65420 $D=1
M196 8 360 1266 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=51530 $D=1
M197 8 361 1267 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=56160 $D=1
M198 8 362 1268 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=60790 $D=1
M199 8 363 1269 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=65420 $D=1
M200 364 1266 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=51530 $D=1
M201 365 1267 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=56160 $D=1
M202 366 1268 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=60790 $D=1
M203 367 1269 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=65420 $D=1
M204 360 352 364 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=51530 $D=1
M205 361 353 365 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=56160 $D=1
M206 362 354 366 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=60790 $D=1
M207 363 355 367 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=65420 $D=1
M208 364 30 320 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=51530 $D=1
M209 365 30 321 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=56160 $D=1
M210 366 30 322 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=60790 $D=1
M211 367 30 323 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=65420 $D=1
M212 328 31 364 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=51530 $D=1
M213 329 31 365 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=56160 $D=1
M214 330 31 366 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=60790 $D=1
M215 331 31 367 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=65420 $D=1
M216 368 31 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=51530 $D=1
M217 369 31 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=56160 $D=1
M218 370 31 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=60790 $D=1
M219 371 31 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=65420 $D=1
M220 8 32 372 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=51530 $D=1
M221 8 32 373 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=56160 $D=1
M222 8 32 374 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=60790 $D=1
M223 8 32 375 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=65420 $D=1
M224 376 33 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=51530 $D=1
M225 377 33 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=56160 $D=1
M226 378 33 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=60790 $D=1
M227 379 33 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=65420 $D=1
M228 380 32 300 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=51530 $D=1
M229 381 32 301 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=56160 $D=1
M230 382 32 302 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=60790 $D=1
M231 383 32 303 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=65420 $D=1
M232 8 380 1270 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=51530 $D=1
M233 8 381 1271 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=56160 $D=1
M234 8 382 1272 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=60790 $D=1
M235 8 383 1273 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=65420 $D=1
M236 384 1270 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=51530 $D=1
M237 385 1271 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=56160 $D=1
M238 386 1272 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=60790 $D=1
M239 387 1273 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=65420 $D=1
M240 380 372 384 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=51530 $D=1
M241 381 373 385 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=56160 $D=1
M242 382 374 386 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=60790 $D=1
M243 383 375 387 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=65420 $D=1
M244 384 33 320 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=51530 $D=1
M245 385 33 321 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=56160 $D=1
M246 386 33 322 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=60790 $D=1
M247 387 33 323 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=65420 $D=1
M248 328 34 384 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=51530 $D=1
M249 329 34 385 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=56160 $D=1
M250 330 34 386 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=60790 $D=1
M251 331 34 387 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=65420 $D=1
M252 388 34 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=51530 $D=1
M253 389 34 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=56160 $D=1
M254 390 34 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=60790 $D=1
M255 391 34 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=65420 $D=1
M256 8 35 392 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=51530 $D=1
M257 8 35 393 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=56160 $D=1
M258 8 35 394 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=60790 $D=1
M259 8 35 395 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=65420 $D=1
M260 396 36 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=51530 $D=1
M261 397 36 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=56160 $D=1
M262 398 36 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=60790 $D=1
M263 399 36 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=65420 $D=1
M264 400 35 300 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=51530 $D=1
M265 401 35 301 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=56160 $D=1
M266 402 35 302 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=60790 $D=1
M267 403 35 303 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=65420 $D=1
M268 8 400 1274 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=51530 $D=1
M269 8 401 1275 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=56160 $D=1
M270 8 402 1276 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=60790 $D=1
M271 8 403 1277 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=65420 $D=1
M272 404 1274 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=51530 $D=1
M273 405 1275 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=56160 $D=1
M274 406 1276 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=60790 $D=1
M275 407 1277 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=65420 $D=1
M276 400 392 404 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=51530 $D=1
M277 401 393 405 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=56160 $D=1
M278 402 394 406 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=60790 $D=1
M279 403 395 407 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=65420 $D=1
M280 404 36 320 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=51530 $D=1
M281 405 36 321 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=56160 $D=1
M282 406 36 322 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=60790 $D=1
M283 407 36 323 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=65420 $D=1
M284 328 37 404 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=51530 $D=1
M285 329 37 405 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=56160 $D=1
M286 330 37 406 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=60790 $D=1
M287 331 37 407 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=65420 $D=1
M288 408 37 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=51530 $D=1
M289 409 37 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=56160 $D=1
M290 410 37 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=60790 $D=1
M291 411 37 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=65420 $D=1
M292 8 38 412 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=51530 $D=1
M293 8 38 413 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=56160 $D=1
M294 8 38 414 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=60790 $D=1
M295 8 38 415 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=65420 $D=1
M296 416 39 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=51530 $D=1
M297 417 39 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=56160 $D=1
M298 418 39 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=60790 $D=1
M299 419 39 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=65420 $D=1
M300 420 38 300 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=51530 $D=1
M301 421 38 301 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=56160 $D=1
M302 422 38 302 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=60790 $D=1
M303 423 38 303 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=65420 $D=1
M304 8 420 1278 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=51530 $D=1
M305 8 421 1279 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=56160 $D=1
M306 8 422 1280 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=60790 $D=1
M307 8 423 1281 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=65420 $D=1
M308 424 1278 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=51530 $D=1
M309 425 1279 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=56160 $D=1
M310 426 1280 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=60790 $D=1
M311 427 1281 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=65420 $D=1
M312 420 412 424 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=51530 $D=1
M313 421 413 425 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=56160 $D=1
M314 422 414 426 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=60790 $D=1
M315 423 415 427 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=65420 $D=1
M316 424 39 320 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=51530 $D=1
M317 425 39 321 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=56160 $D=1
M318 426 39 322 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=60790 $D=1
M319 427 39 323 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=65420 $D=1
M320 328 40 424 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=51530 $D=1
M321 329 40 425 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=56160 $D=1
M322 330 40 426 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=60790 $D=1
M323 331 40 427 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=65420 $D=1
M324 428 40 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=51530 $D=1
M325 429 40 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=56160 $D=1
M326 430 40 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=60790 $D=1
M327 431 40 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=65420 $D=1
M328 8 41 432 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=51530 $D=1
M329 8 41 433 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=56160 $D=1
M330 8 41 434 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=60790 $D=1
M331 8 41 435 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=65420 $D=1
M332 436 42 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=51530 $D=1
M333 437 42 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=56160 $D=1
M334 438 42 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=60790 $D=1
M335 439 42 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=65420 $D=1
M336 440 41 300 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=51530 $D=1
M337 441 41 301 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=56160 $D=1
M338 442 41 302 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=60790 $D=1
M339 443 41 303 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=65420 $D=1
M340 8 440 1282 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=51530 $D=1
M341 8 441 1283 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=56160 $D=1
M342 8 442 1284 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=60790 $D=1
M343 8 443 1285 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=65420 $D=1
M344 444 1282 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=51530 $D=1
M345 445 1283 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=56160 $D=1
M346 446 1284 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=60790 $D=1
M347 447 1285 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=65420 $D=1
M348 440 432 444 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=51530 $D=1
M349 441 433 445 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=56160 $D=1
M350 442 434 446 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=60790 $D=1
M351 443 435 447 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=65420 $D=1
M352 444 42 320 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=51530 $D=1
M353 445 42 321 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=56160 $D=1
M354 446 42 322 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=60790 $D=1
M355 447 42 323 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=65420 $D=1
M356 328 43 444 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=51530 $D=1
M357 329 43 445 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=56160 $D=1
M358 330 43 446 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=60790 $D=1
M359 331 43 447 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=65420 $D=1
M360 448 43 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=51530 $D=1
M361 449 43 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=56160 $D=1
M362 450 43 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=60790 $D=1
M363 451 43 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=65420 $D=1
M364 8 44 452 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=51530 $D=1
M365 8 44 453 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=56160 $D=1
M366 8 44 454 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=60790 $D=1
M367 8 44 455 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=65420 $D=1
M368 456 45 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=51530 $D=1
M369 457 45 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=56160 $D=1
M370 458 45 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=60790 $D=1
M371 459 45 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=65420 $D=1
M372 460 44 300 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=51530 $D=1
M373 461 44 301 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=56160 $D=1
M374 462 44 302 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=60790 $D=1
M375 463 44 303 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=65420 $D=1
M376 8 460 1286 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=51530 $D=1
M377 8 461 1287 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=56160 $D=1
M378 8 462 1288 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=60790 $D=1
M379 8 463 1289 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=65420 $D=1
M380 464 1286 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=51530 $D=1
M381 465 1287 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=56160 $D=1
M382 466 1288 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=60790 $D=1
M383 467 1289 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=65420 $D=1
M384 460 452 464 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=51530 $D=1
M385 461 453 465 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=56160 $D=1
M386 462 454 466 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=60790 $D=1
M387 463 455 467 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=65420 $D=1
M388 464 45 320 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=51530 $D=1
M389 465 45 321 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=56160 $D=1
M390 466 45 322 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=60790 $D=1
M391 467 45 323 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=65420 $D=1
M392 328 46 464 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=51530 $D=1
M393 329 46 465 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=56160 $D=1
M394 330 46 466 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=60790 $D=1
M395 331 46 467 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=65420 $D=1
M396 468 46 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=51530 $D=1
M397 469 46 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=56160 $D=1
M398 470 46 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=60790 $D=1
M399 471 46 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=65420 $D=1
M400 8 47 472 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=51530 $D=1
M401 8 47 473 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=56160 $D=1
M402 8 47 474 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=60790 $D=1
M403 8 47 475 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=65420 $D=1
M404 476 48 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=51530 $D=1
M405 477 48 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=56160 $D=1
M406 478 48 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=60790 $D=1
M407 479 48 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=65420 $D=1
M408 480 47 300 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=51530 $D=1
M409 481 47 301 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=56160 $D=1
M410 482 47 302 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=60790 $D=1
M411 483 47 303 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=65420 $D=1
M412 8 480 1290 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=51530 $D=1
M413 8 481 1291 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=56160 $D=1
M414 8 482 1292 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=60790 $D=1
M415 8 483 1293 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=65420 $D=1
M416 484 1290 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=51530 $D=1
M417 485 1291 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=56160 $D=1
M418 486 1292 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=60790 $D=1
M419 487 1293 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=65420 $D=1
M420 480 472 484 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=51530 $D=1
M421 481 473 485 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=56160 $D=1
M422 482 474 486 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=60790 $D=1
M423 483 475 487 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=65420 $D=1
M424 484 48 320 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=51530 $D=1
M425 485 48 321 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=56160 $D=1
M426 486 48 322 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=60790 $D=1
M427 487 48 323 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=65420 $D=1
M428 328 49 484 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=51530 $D=1
M429 329 49 485 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=56160 $D=1
M430 330 49 486 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=60790 $D=1
M431 331 49 487 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=65420 $D=1
M432 488 49 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=51530 $D=1
M433 489 49 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=56160 $D=1
M434 490 49 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=60790 $D=1
M435 491 49 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=65420 $D=1
M436 8 50 492 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=51530 $D=1
M437 8 50 493 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=56160 $D=1
M438 8 50 494 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=60790 $D=1
M439 8 50 495 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=65420 $D=1
M440 496 51 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=51530 $D=1
M441 497 51 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=56160 $D=1
M442 498 51 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=60790 $D=1
M443 499 51 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=65420 $D=1
M444 500 50 300 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=51530 $D=1
M445 501 50 301 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=56160 $D=1
M446 502 50 302 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=60790 $D=1
M447 503 50 303 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=65420 $D=1
M448 8 500 1294 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=51530 $D=1
M449 8 501 1295 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=56160 $D=1
M450 8 502 1296 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=60790 $D=1
M451 8 503 1297 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=65420 $D=1
M452 504 1294 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=51530 $D=1
M453 505 1295 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=56160 $D=1
M454 506 1296 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=60790 $D=1
M455 507 1297 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=65420 $D=1
M456 500 492 504 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=51530 $D=1
M457 501 493 505 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=56160 $D=1
M458 502 494 506 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=60790 $D=1
M459 503 495 507 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=65420 $D=1
M460 504 51 320 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=51530 $D=1
M461 505 51 321 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=56160 $D=1
M462 506 51 322 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=60790 $D=1
M463 507 51 323 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=65420 $D=1
M464 328 52 504 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=51530 $D=1
M465 329 52 505 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=56160 $D=1
M466 330 52 506 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=60790 $D=1
M467 331 52 507 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=65420 $D=1
M468 508 52 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=51530 $D=1
M469 509 52 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=56160 $D=1
M470 510 52 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=60790 $D=1
M471 511 52 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=65420 $D=1
M472 8 53 512 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=51530 $D=1
M473 8 53 513 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=56160 $D=1
M474 8 53 514 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=60790 $D=1
M475 8 53 515 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=65420 $D=1
M476 516 54 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=51530 $D=1
M477 517 54 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=56160 $D=1
M478 518 54 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=60790 $D=1
M479 519 54 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=65420 $D=1
M480 520 53 300 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=51530 $D=1
M481 521 53 301 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=56160 $D=1
M482 522 53 302 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=60790 $D=1
M483 523 53 303 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=65420 $D=1
M484 8 520 1298 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=51530 $D=1
M485 8 521 1299 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=56160 $D=1
M486 8 522 1300 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=60790 $D=1
M487 8 523 1301 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=65420 $D=1
M488 524 1298 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=51530 $D=1
M489 525 1299 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=56160 $D=1
M490 526 1300 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=60790 $D=1
M491 527 1301 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=65420 $D=1
M492 520 512 524 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=51530 $D=1
M493 521 513 525 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=56160 $D=1
M494 522 514 526 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=60790 $D=1
M495 523 515 527 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=65420 $D=1
M496 524 54 320 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=51530 $D=1
M497 525 54 321 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=56160 $D=1
M498 526 54 322 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=60790 $D=1
M499 527 54 323 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=65420 $D=1
M500 328 55 524 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=51530 $D=1
M501 329 55 525 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=56160 $D=1
M502 330 55 526 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=60790 $D=1
M503 331 55 527 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=65420 $D=1
M504 528 55 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=51530 $D=1
M505 529 55 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=56160 $D=1
M506 530 55 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=60790 $D=1
M507 531 55 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=65420 $D=1
M508 8 56 532 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=51530 $D=1
M509 8 56 533 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=56160 $D=1
M510 8 56 534 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=60790 $D=1
M511 8 56 535 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=65420 $D=1
M512 536 57 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=51530 $D=1
M513 537 57 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=56160 $D=1
M514 538 57 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=60790 $D=1
M515 539 57 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=65420 $D=1
M516 540 56 300 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=51530 $D=1
M517 541 56 301 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=56160 $D=1
M518 542 56 302 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=60790 $D=1
M519 543 56 303 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=65420 $D=1
M520 8 540 1302 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=51530 $D=1
M521 8 541 1303 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=56160 $D=1
M522 8 542 1304 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=60790 $D=1
M523 8 543 1305 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=65420 $D=1
M524 544 1302 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=51530 $D=1
M525 545 1303 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=56160 $D=1
M526 546 1304 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=60790 $D=1
M527 547 1305 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=65420 $D=1
M528 540 532 544 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=51530 $D=1
M529 541 533 545 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=56160 $D=1
M530 542 534 546 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=60790 $D=1
M531 543 535 547 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=65420 $D=1
M532 544 57 320 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=51530 $D=1
M533 545 57 321 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=56160 $D=1
M534 546 57 322 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=60790 $D=1
M535 547 57 323 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=65420 $D=1
M536 328 58 544 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=51530 $D=1
M537 329 58 545 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=56160 $D=1
M538 330 58 546 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=60790 $D=1
M539 331 58 547 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=65420 $D=1
M540 548 58 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=51530 $D=1
M541 549 58 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=56160 $D=1
M542 550 58 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=60790 $D=1
M543 551 58 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=65420 $D=1
M544 8 59 552 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=51530 $D=1
M545 8 59 553 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=56160 $D=1
M546 8 59 554 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=60790 $D=1
M547 8 59 555 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=65420 $D=1
M548 556 60 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=51530 $D=1
M549 557 60 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=56160 $D=1
M550 558 60 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=60790 $D=1
M551 559 60 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=65420 $D=1
M552 560 59 300 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=51530 $D=1
M553 561 59 301 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=56160 $D=1
M554 562 59 302 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=60790 $D=1
M555 563 59 303 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=65420 $D=1
M556 8 560 1306 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=51530 $D=1
M557 8 561 1307 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=56160 $D=1
M558 8 562 1308 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=60790 $D=1
M559 8 563 1309 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=65420 $D=1
M560 564 1306 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=51530 $D=1
M561 565 1307 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=56160 $D=1
M562 566 1308 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=60790 $D=1
M563 567 1309 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=65420 $D=1
M564 560 552 564 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=51530 $D=1
M565 561 553 565 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=56160 $D=1
M566 562 554 566 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=60790 $D=1
M567 563 555 567 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=65420 $D=1
M568 564 60 320 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=51530 $D=1
M569 565 60 321 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=56160 $D=1
M570 566 60 322 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=60790 $D=1
M571 567 60 323 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=65420 $D=1
M572 328 61 564 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=51530 $D=1
M573 329 61 565 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=56160 $D=1
M574 330 61 566 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=60790 $D=1
M575 331 61 567 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=65420 $D=1
M576 568 61 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=51530 $D=1
M577 569 61 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=56160 $D=1
M578 570 61 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=60790 $D=1
M579 571 61 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=65420 $D=1
M580 8 62 572 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=51530 $D=1
M581 8 62 573 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=56160 $D=1
M582 8 62 574 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=60790 $D=1
M583 8 62 575 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=65420 $D=1
M584 576 63 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=51530 $D=1
M585 577 63 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=56160 $D=1
M586 578 63 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=60790 $D=1
M587 579 63 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=65420 $D=1
M588 580 62 300 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=51530 $D=1
M589 581 62 301 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=56160 $D=1
M590 582 62 302 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=60790 $D=1
M591 583 62 303 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=65420 $D=1
M592 8 580 1310 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=51530 $D=1
M593 8 581 1311 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=56160 $D=1
M594 8 582 1312 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=60790 $D=1
M595 8 583 1313 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=65420 $D=1
M596 584 1310 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=51530 $D=1
M597 585 1311 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=56160 $D=1
M598 586 1312 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=60790 $D=1
M599 587 1313 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=65420 $D=1
M600 580 572 584 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=51530 $D=1
M601 581 573 585 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=56160 $D=1
M602 582 574 586 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=60790 $D=1
M603 583 575 587 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=65420 $D=1
M604 584 63 320 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=51530 $D=1
M605 585 63 321 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=56160 $D=1
M606 586 63 322 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=60790 $D=1
M607 587 63 323 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=65420 $D=1
M608 328 64 584 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=51530 $D=1
M609 329 64 585 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=56160 $D=1
M610 330 64 586 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=60790 $D=1
M611 331 64 587 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=65420 $D=1
M612 588 64 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=51530 $D=1
M613 589 64 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=56160 $D=1
M614 590 64 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=60790 $D=1
M615 591 64 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=65420 $D=1
M616 8 65 592 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=51530 $D=1
M617 8 65 593 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=56160 $D=1
M618 8 65 594 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=60790 $D=1
M619 8 65 595 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=65420 $D=1
M620 596 66 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=51530 $D=1
M621 597 66 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=56160 $D=1
M622 598 66 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=60790 $D=1
M623 599 66 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=65420 $D=1
M624 600 65 300 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=51530 $D=1
M625 601 65 301 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=56160 $D=1
M626 602 65 302 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=60790 $D=1
M627 603 65 303 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=65420 $D=1
M628 8 600 1314 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=51530 $D=1
M629 8 601 1315 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=56160 $D=1
M630 8 602 1316 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=60790 $D=1
M631 8 603 1317 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=65420 $D=1
M632 604 1314 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=51530 $D=1
M633 605 1315 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=56160 $D=1
M634 606 1316 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=60790 $D=1
M635 607 1317 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=65420 $D=1
M636 600 592 604 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=51530 $D=1
M637 601 593 605 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=56160 $D=1
M638 602 594 606 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=60790 $D=1
M639 603 595 607 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=65420 $D=1
M640 604 66 320 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=51530 $D=1
M641 605 66 321 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=56160 $D=1
M642 606 66 322 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=60790 $D=1
M643 607 66 323 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=65420 $D=1
M644 328 67 604 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=51530 $D=1
M645 329 67 605 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=56160 $D=1
M646 330 67 606 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=60790 $D=1
M647 331 67 607 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=65420 $D=1
M648 608 67 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=51530 $D=1
M649 609 67 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=56160 $D=1
M650 610 67 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=60790 $D=1
M651 611 67 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=65420 $D=1
M652 8 68 612 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=51530 $D=1
M653 8 68 613 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=56160 $D=1
M654 8 68 614 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=60790 $D=1
M655 8 68 615 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=65420 $D=1
M656 616 69 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=51530 $D=1
M657 617 69 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=56160 $D=1
M658 618 69 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=60790 $D=1
M659 619 69 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=65420 $D=1
M660 620 68 300 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=51530 $D=1
M661 621 68 301 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=56160 $D=1
M662 622 68 302 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=60790 $D=1
M663 623 68 303 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=65420 $D=1
M664 8 620 1318 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=51530 $D=1
M665 8 621 1319 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=56160 $D=1
M666 8 622 1320 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=60790 $D=1
M667 8 623 1321 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=65420 $D=1
M668 624 1318 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=51530 $D=1
M669 625 1319 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=56160 $D=1
M670 626 1320 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=60790 $D=1
M671 627 1321 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=65420 $D=1
M672 620 612 624 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=51530 $D=1
M673 621 613 625 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=56160 $D=1
M674 622 614 626 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=60790 $D=1
M675 623 615 627 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=65420 $D=1
M676 624 69 320 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=51530 $D=1
M677 625 69 321 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=56160 $D=1
M678 626 69 322 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=60790 $D=1
M679 627 69 323 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=65420 $D=1
M680 328 70 624 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=51530 $D=1
M681 329 70 625 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=56160 $D=1
M682 330 70 626 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=60790 $D=1
M683 331 70 627 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=65420 $D=1
M684 628 70 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=51530 $D=1
M685 629 70 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=56160 $D=1
M686 630 70 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=60790 $D=1
M687 631 70 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=65420 $D=1
M688 8 71 632 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=51530 $D=1
M689 8 71 633 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=56160 $D=1
M690 8 71 634 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=60790 $D=1
M691 8 71 635 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=65420 $D=1
M692 636 72 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=51530 $D=1
M693 637 72 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=56160 $D=1
M694 638 72 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=60790 $D=1
M695 639 72 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=65420 $D=1
M696 640 71 300 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=51530 $D=1
M697 641 71 301 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=56160 $D=1
M698 642 71 302 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=60790 $D=1
M699 643 71 303 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=65420 $D=1
M700 8 640 1322 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=51530 $D=1
M701 8 641 1323 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=56160 $D=1
M702 8 642 1324 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=60790 $D=1
M703 8 643 1325 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=65420 $D=1
M704 644 1322 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=51530 $D=1
M705 645 1323 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=56160 $D=1
M706 646 1324 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=60790 $D=1
M707 647 1325 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=65420 $D=1
M708 640 632 644 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=51530 $D=1
M709 641 633 645 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=56160 $D=1
M710 642 634 646 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=60790 $D=1
M711 643 635 647 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=65420 $D=1
M712 644 72 320 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=51530 $D=1
M713 645 72 321 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=56160 $D=1
M714 646 72 322 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=60790 $D=1
M715 647 72 323 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=65420 $D=1
M716 328 73 644 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=51530 $D=1
M717 329 73 645 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=56160 $D=1
M718 330 73 646 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=60790 $D=1
M719 331 73 647 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=65420 $D=1
M720 648 73 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=51530 $D=1
M721 649 73 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=56160 $D=1
M722 650 73 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=60790 $D=1
M723 651 73 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=65420 $D=1
M724 8 74 652 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=51530 $D=1
M725 8 74 653 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=56160 $D=1
M726 8 74 654 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=60790 $D=1
M727 8 74 655 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=65420 $D=1
M728 656 75 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=51530 $D=1
M729 657 75 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=56160 $D=1
M730 658 75 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=60790 $D=1
M731 659 75 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=65420 $D=1
M732 660 74 300 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=51530 $D=1
M733 661 74 301 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=56160 $D=1
M734 662 74 302 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=60790 $D=1
M735 663 74 303 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=65420 $D=1
M736 8 660 1326 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=51530 $D=1
M737 8 661 1327 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=56160 $D=1
M738 8 662 1328 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=60790 $D=1
M739 8 663 1329 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=65420 $D=1
M740 664 1326 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=51530 $D=1
M741 665 1327 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=56160 $D=1
M742 666 1328 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=60790 $D=1
M743 667 1329 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=65420 $D=1
M744 660 652 664 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=51530 $D=1
M745 661 653 665 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=56160 $D=1
M746 662 654 666 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=60790 $D=1
M747 663 655 667 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=65420 $D=1
M748 664 75 320 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=51530 $D=1
M749 665 75 321 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=56160 $D=1
M750 666 75 322 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=60790 $D=1
M751 667 75 323 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=65420 $D=1
M752 328 76 664 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=51530 $D=1
M753 329 76 665 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=56160 $D=1
M754 330 76 666 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=60790 $D=1
M755 331 76 667 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=65420 $D=1
M756 668 76 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=51530 $D=1
M757 669 76 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=56160 $D=1
M758 670 76 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=60790 $D=1
M759 671 76 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=65420 $D=1
M760 8 77 672 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=51530 $D=1
M761 8 77 673 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=56160 $D=1
M762 8 77 674 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=60790 $D=1
M763 8 77 675 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=65420 $D=1
M764 676 78 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=51530 $D=1
M765 677 78 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=56160 $D=1
M766 678 78 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=60790 $D=1
M767 679 78 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=65420 $D=1
M768 680 77 300 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=51530 $D=1
M769 681 77 301 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=56160 $D=1
M770 682 77 302 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=60790 $D=1
M771 683 77 303 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=65420 $D=1
M772 8 680 1330 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=51530 $D=1
M773 8 681 1331 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=56160 $D=1
M774 8 682 1332 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=60790 $D=1
M775 8 683 1333 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=65420 $D=1
M776 684 1330 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=51530 $D=1
M777 685 1331 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=56160 $D=1
M778 686 1332 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=60790 $D=1
M779 687 1333 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=65420 $D=1
M780 680 672 684 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=51530 $D=1
M781 681 673 685 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=56160 $D=1
M782 682 674 686 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=60790 $D=1
M783 683 675 687 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=65420 $D=1
M784 684 78 320 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=51530 $D=1
M785 685 78 321 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=56160 $D=1
M786 686 78 322 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=60790 $D=1
M787 687 78 323 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=65420 $D=1
M788 328 79 684 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=51530 $D=1
M789 329 79 685 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=56160 $D=1
M790 330 79 686 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=60790 $D=1
M791 331 79 687 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=65420 $D=1
M792 688 79 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=51530 $D=1
M793 689 79 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=56160 $D=1
M794 690 79 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=60790 $D=1
M795 691 79 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=65420 $D=1
M796 8 80 692 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=51530 $D=1
M797 8 80 693 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=56160 $D=1
M798 8 80 694 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=60790 $D=1
M799 8 80 695 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=65420 $D=1
M800 696 81 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=51530 $D=1
M801 697 81 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=56160 $D=1
M802 698 81 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=60790 $D=1
M803 699 81 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=65420 $D=1
M804 700 80 300 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=51530 $D=1
M805 701 80 301 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=56160 $D=1
M806 702 80 302 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=60790 $D=1
M807 703 80 303 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=65420 $D=1
M808 8 700 1334 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=51530 $D=1
M809 8 701 1335 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=56160 $D=1
M810 8 702 1336 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=60790 $D=1
M811 8 703 1337 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=65420 $D=1
M812 704 1334 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=51530 $D=1
M813 705 1335 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=56160 $D=1
M814 706 1336 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=60790 $D=1
M815 707 1337 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=65420 $D=1
M816 700 692 704 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=51530 $D=1
M817 701 693 705 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=56160 $D=1
M818 702 694 706 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=60790 $D=1
M819 703 695 707 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=65420 $D=1
M820 704 81 320 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=51530 $D=1
M821 705 81 321 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=56160 $D=1
M822 706 81 322 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=60790 $D=1
M823 707 81 323 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=65420 $D=1
M824 328 82 704 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=51530 $D=1
M825 329 82 705 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=56160 $D=1
M826 330 82 706 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=60790 $D=1
M827 331 82 707 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=65420 $D=1
M828 708 82 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=51530 $D=1
M829 709 82 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=56160 $D=1
M830 710 82 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=60790 $D=1
M831 711 82 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=65420 $D=1
M832 8 83 712 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=51530 $D=1
M833 8 83 713 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=56160 $D=1
M834 8 83 714 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=60790 $D=1
M835 8 83 715 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=65420 $D=1
M836 716 84 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=51530 $D=1
M837 717 84 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=56160 $D=1
M838 718 84 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=60790 $D=1
M839 719 84 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=65420 $D=1
M840 720 83 300 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=51530 $D=1
M841 721 83 301 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=56160 $D=1
M842 722 83 302 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=60790 $D=1
M843 723 83 303 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=65420 $D=1
M844 8 720 1338 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=51530 $D=1
M845 8 721 1339 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=56160 $D=1
M846 8 722 1340 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=60790 $D=1
M847 8 723 1341 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=65420 $D=1
M848 724 1338 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=51530 $D=1
M849 725 1339 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=56160 $D=1
M850 726 1340 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=60790 $D=1
M851 727 1341 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=65420 $D=1
M852 720 712 724 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=51530 $D=1
M853 721 713 725 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=56160 $D=1
M854 722 714 726 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=60790 $D=1
M855 723 715 727 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=65420 $D=1
M856 724 84 320 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=51530 $D=1
M857 725 84 321 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=56160 $D=1
M858 726 84 322 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=60790 $D=1
M859 727 84 323 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=65420 $D=1
M860 328 85 724 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=51530 $D=1
M861 329 85 725 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=56160 $D=1
M862 330 85 726 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=60790 $D=1
M863 331 85 727 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=65420 $D=1
M864 728 85 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=51530 $D=1
M865 729 85 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=56160 $D=1
M866 730 85 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=60790 $D=1
M867 731 85 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=65420 $D=1
M868 8 86 732 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=51530 $D=1
M869 8 86 733 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=56160 $D=1
M870 8 86 734 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=60790 $D=1
M871 8 86 735 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=65420 $D=1
M872 736 87 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=51530 $D=1
M873 737 87 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=56160 $D=1
M874 738 87 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=60790 $D=1
M875 739 87 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=65420 $D=1
M876 740 86 300 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=51530 $D=1
M877 741 86 301 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=56160 $D=1
M878 742 86 302 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=60790 $D=1
M879 743 86 303 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=65420 $D=1
M880 8 740 1342 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=51530 $D=1
M881 8 741 1343 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=56160 $D=1
M882 8 742 1344 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=60790 $D=1
M883 8 743 1345 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=65420 $D=1
M884 744 1342 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=51530 $D=1
M885 745 1343 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=56160 $D=1
M886 746 1344 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=60790 $D=1
M887 747 1345 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=65420 $D=1
M888 740 732 744 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=51530 $D=1
M889 741 733 745 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=56160 $D=1
M890 742 734 746 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=60790 $D=1
M891 743 735 747 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=65420 $D=1
M892 744 87 320 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=51530 $D=1
M893 745 87 321 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=56160 $D=1
M894 746 87 322 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=60790 $D=1
M895 747 87 323 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=65420 $D=1
M896 328 88 744 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=51530 $D=1
M897 329 88 745 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=56160 $D=1
M898 330 88 746 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=60790 $D=1
M899 331 88 747 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=65420 $D=1
M900 748 88 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=51530 $D=1
M901 749 88 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=56160 $D=1
M902 750 88 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=60790 $D=1
M903 751 88 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=65420 $D=1
M904 8 89 752 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=51530 $D=1
M905 8 89 753 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=56160 $D=1
M906 8 89 754 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=60790 $D=1
M907 8 89 755 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=65420 $D=1
M908 756 90 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=51530 $D=1
M909 757 90 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=56160 $D=1
M910 758 90 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=60790 $D=1
M911 759 90 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=65420 $D=1
M912 760 89 300 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=51530 $D=1
M913 761 89 301 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=56160 $D=1
M914 762 89 302 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=60790 $D=1
M915 763 89 303 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=65420 $D=1
M916 8 760 1346 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=51530 $D=1
M917 8 761 1347 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=56160 $D=1
M918 8 762 1348 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=60790 $D=1
M919 8 763 1349 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=65420 $D=1
M920 764 1346 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=51530 $D=1
M921 765 1347 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=56160 $D=1
M922 766 1348 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=60790 $D=1
M923 767 1349 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=65420 $D=1
M924 760 752 764 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=51530 $D=1
M925 761 753 765 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=56160 $D=1
M926 762 754 766 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=60790 $D=1
M927 763 755 767 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=65420 $D=1
M928 764 90 320 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=51530 $D=1
M929 765 90 321 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=56160 $D=1
M930 766 90 322 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=60790 $D=1
M931 767 90 323 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=65420 $D=1
M932 328 91 764 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=51530 $D=1
M933 329 91 765 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=56160 $D=1
M934 330 91 766 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=60790 $D=1
M935 331 91 767 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=65420 $D=1
M936 768 91 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=51530 $D=1
M937 769 91 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=56160 $D=1
M938 770 91 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=60790 $D=1
M939 771 91 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=65420 $D=1
M940 8 92 772 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=51530 $D=1
M941 8 92 773 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=56160 $D=1
M942 8 92 774 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=60790 $D=1
M943 8 92 775 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=65420 $D=1
M944 776 93 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=51530 $D=1
M945 777 93 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=56160 $D=1
M946 778 93 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=60790 $D=1
M947 779 93 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=65420 $D=1
M948 780 92 300 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=51530 $D=1
M949 781 92 301 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=56160 $D=1
M950 782 92 302 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=60790 $D=1
M951 783 92 303 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=65420 $D=1
M952 8 780 1350 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=51530 $D=1
M953 8 781 1351 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=56160 $D=1
M954 8 782 1352 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=60790 $D=1
M955 8 783 1353 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=65420 $D=1
M956 784 1350 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=51530 $D=1
M957 785 1351 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=56160 $D=1
M958 786 1352 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=60790 $D=1
M959 787 1353 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=65420 $D=1
M960 780 772 784 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=51530 $D=1
M961 781 773 785 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=56160 $D=1
M962 782 774 786 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=60790 $D=1
M963 783 775 787 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=65420 $D=1
M964 784 93 320 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=51530 $D=1
M965 785 93 321 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=56160 $D=1
M966 786 93 322 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=60790 $D=1
M967 787 93 323 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=65420 $D=1
M968 328 94 784 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=51530 $D=1
M969 329 94 785 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=56160 $D=1
M970 330 94 786 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=60790 $D=1
M971 331 94 787 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=65420 $D=1
M972 788 94 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=51530 $D=1
M973 789 94 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=56160 $D=1
M974 790 94 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=60790 $D=1
M975 791 94 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=65420 $D=1
M976 8 95 792 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=51530 $D=1
M977 8 95 793 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=56160 $D=1
M978 8 95 794 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=60790 $D=1
M979 8 95 795 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=65420 $D=1
M980 796 96 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=51530 $D=1
M981 797 96 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=56160 $D=1
M982 798 96 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=60790 $D=1
M983 799 96 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=65420 $D=1
M984 800 95 300 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=51530 $D=1
M985 801 95 301 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=56160 $D=1
M986 802 95 302 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=60790 $D=1
M987 803 95 303 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=65420 $D=1
M988 8 800 1354 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=51530 $D=1
M989 8 801 1355 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=56160 $D=1
M990 8 802 1356 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=60790 $D=1
M991 8 803 1357 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=65420 $D=1
M992 804 1354 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=51530 $D=1
M993 805 1355 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=56160 $D=1
M994 806 1356 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=60790 $D=1
M995 807 1357 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=65420 $D=1
M996 800 792 804 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=51530 $D=1
M997 801 793 805 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=56160 $D=1
M998 802 794 806 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=60790 $D=1
M999 803 795 807 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=65420 $D=1
M1000 804 96 320 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=51530 $D=1
M1001 805 96 321 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=56160 $D=1
M1002 806 96 322 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=60790 $D=1
M1003 807 96 323 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=65420 $D=1
M1004 328 97 804 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=51530 $D=1
M1005 329 97 805 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=56160 $D=1
M1006 330 97 806 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=60790 $D=1
M1007 331 97 807 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=65420 $D=1
M1008 808 97 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=51530 $D=1
M1009 809 97 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=56160 $D=1
M1010 810 97 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=60790 $D=1
M1011 811 97 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=65420 $D=1
M1012 8 98 812 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=51530 $D=1
M1013 8 98 813 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=56160 $D=1
M1014 8 98 814 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=60790 $D=1
M1015 8 98 815 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=65420 $D=1
M1016 816 99 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=51530 $D=1
M1017 817 99 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=56160 $D=1
M1018 818 99 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=60790 $D=1
M1019 819 99 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=65420 $D=1
M1020 820 98 300 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=51530 $D=1
M1021 821 98 301 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=56160 $D=1
M1022 822 98 302 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=60790 $D=1
M1023 823 98 303 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=65420 $D=1
M1024 8 820 1358 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=51530 $D=1
M1025 8 821 1359 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=56160 $D=1
M1026 8 822 1360 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=60790 $D=1
M1027 8 823 1361 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=65420 $D=1
M1028 824 1358 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=51530 $D=1
M1029 825 1359 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=56160 $D=1
M1030 826 1360 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=60790 $D=1
M1031 827 1361 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=65420 $D=1
M1032 820 812 824 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=51530 $D=1
M1033 821 813 825 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=56160 $D=1
M1034 822 814 826 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=60790 $D=1
M1035 823 815 827 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=65420 $D=1
M1036 824 99 320 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=51530 $D=1
M1037 825 99 321 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=56160 $D=1
M1038 826 99 322 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=60790 $D=1
M1039 827 99 323 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=65420 $D=1
M1040 328 100 824 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=51530 $D=1
M1041 329 100 825 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=56160 $D=1
M1042 330 100 826 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=60790 $D=1
M1043 331 100 827 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=65420 $D=1
M1044 828 100 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=51530 $D=1
M1045 829 100 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=56160 $D=1
M1046 830 100 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=60790 $D=1
M1047 831 100 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=65420 $D=1
M1048 8 101 832 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=51530 $D=1
M1049 8 101 833 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=56160 $D=1
M1050 8 101 834 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=60790 $D=1
M1051 8 101 835 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=65420 $D=1
M1052 836 102 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=51530 $D=1
M1053 837 102 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=56160 $D=1
M1054 838 102 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=60790 $D=1
M1055 839 102 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=65420 $D=1
M1056 840 101 300 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=51530 $D=1
M1057 841 101 301 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=56160 $D=1
M1058 842 101 302 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=60790 $D=1
M1059 843 101 303 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=65420 $D=1
M1060 8 840 1362 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=51530 $D=1
M1061 8 841 1363 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=56160 $D=1
M1062 8 842 1364 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=60790 $D=1
M1063 8 843 1365 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=65420 $D=1
M1064 844 1362 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=51530 $D=1
M1065 845 1363 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=56160 $D=1
M1066 846 1364 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=60790 $D=1
M1067 847 1365 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=65420 $D=1
M1068 840 832 844 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=51530 $D=1
M1069 841 833 845 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=56160 $D=1
M1070 842 834 846 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=60790 $D=1
M1071 843 835 847 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=65420 $D=1
M1072 844 102 320 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=51530 $D=1
M1073 845 102 321 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=56160 $D=1
M1074 846 102 322 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=60790 $D=1
M1075 847 102 323 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=65420 $D=1
M1076 328 103 844 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=51530 $D=1
M1077 329 103 845 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=56160 $D=1
M1078 330 103 846 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=60790 $D=1
M1079 331 103 847 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=65420 $D=1
M1080 848 103 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=51530 $D=1
M1081 849 103 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=56160 $D=1
M1082 850 103 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=60790 $D=1
M1083 851 103 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=65420 $D=1
M1084 8 104 852 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=51530 $D=1
M1085 8 104 853 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=56160 $D=1
M1086 8 104 854 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=60790 $D=1
M1087 8 104 855 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=65420 $D=1
M1088 856 105 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=51530 $D=1
M1089 857 105 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=56160 $D=1
M1090 858 105 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=60790 $D=1
M1091 859 105 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=65420 $D=1
M1092 860 104 300 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=51530 $D=1
M1093 861 104 301 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=56160 $D=1
M1094 862 104 302 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=60790 $D=1
M1095 863 104 303 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=65420 $D=1
M1096 8 860 1366 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=51530 $D=1
M1097 8 861 1367 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=56160 $D=1
M1098 8 862 1368 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=60790 $D=1
M1099 8 863 1369 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=65420 $D=1
M1100 864 1366 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=51530 $D=1
M1101 865 1367 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=56160 $D=1
M1102 866 1368 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=60790 $D=1
M1103 867 1369 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=65420 $D=1
M1104 860 852 864 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=51530 $D=1
M1105 861 853 865 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=56160 $D=1
M1106 862 854 866 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=60790 $D=1
M1107 863 855 867 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=65420 $D=1
M1108 864 105 320 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=51530 $D=1
M1109 865 105 321 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=56160 $D=1
M1110 866 105 322 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=60790 $D=1
M1111 867 105 323 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=65420 $D=1
M1112 328 106 864 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=51530 $D=1
M1113 329 106 865 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=56160 $D=1
M1114 330 106 866 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=60790 $D=1
M1115 331 106 867 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=65420 $D=1
M1116 868 106 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=51530 $D=1
M1117 869 106 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=56160 $D=1
M1118 870 106 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=60790 $D=1
M1119 871 106 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=65420 $D=1
M1120 8 107 872 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=51530 $D=1
M1121 8 107 873 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=56160 $D=1
M1122 8 107 874 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=60790 $D=1
M1123 8 107 875 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=65420 $D=1
M1124 876 108 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=51530 $D=1
M1125 877 108 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=56160 $D=1
M1126 878 108 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=60790 $D=1
M1127 879 108 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=65420 $D=1
M1128 880 107 300 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=51530 $D=1
M1129 881 107 301 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=56160 $D=1
M1130 882 107 302 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=60790 $D=1
M1131 883 107 303 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=65420 $D=1
M1132 8 880 1370 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=51530 $D=1
M1133 8 881 1371 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=56160 $D=1
M1134 8 882 1372 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=60790 $D=1
M1135 8 883 1373 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=65420 $D=1
M1136 884 1370 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=51530 $D=1
M1137 885 1371 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=56160 $D=1
M1138 886 1372 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=60790 $D=1
M1139 887 1373 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=65420 $D=1
M1140 880 872 884 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=51530 $D=1
M1141 881 873 885 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=56160 $D=1
M1142 882 874 886 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=60790 $D=1
M1143 883 875 887 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=65420 $D=1
M1144 884 108 320 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=51530 $D=1
M1145 885 108 321 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=56160 $D=1
M1146 886 108 322 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=60790 $D=1
M1147 887 108 323 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=65420 $D=1
M1148 328 109 884 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=51530 $D=1
M1149 329 109 885 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=56160 $D=1
M1150 330 109 886 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=60790 $D=1
M1151 331 109 887 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=65420 $D=1
M1152 888 109 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=51530 $D=1
M1153 889 109 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=56160 $D=1
M1154 890 109 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=60790 $D=1
M1155 891 109 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=65420 $D=1
M1156 8 110 892 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=51530 $D=1
M1157 8 110 893 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=56160 $D=1
M1158 8 110 894 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=60790 $D=1
M1159 8 110 895 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=65420 $D=1
M1160 896 111 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=51530 $D=1
M1161 897 111 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=56160 $D=1
M1162 898 111 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=60790 $D=1
M1163 899 111 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=65420 $D=1
M1164 900 110 300 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=51530 $D=1
M1165 901 110 301 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=56160 $D=1
M1166 902 110 302 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=60790 $D=1
M1167 903 110 303 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=65420 $D=1
M1168 8 900 1374 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=51530 $D=1
M1169 8 901 1375 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=56160 $D=1
M1170 8 902 1376 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=60790 $D=1
M1171 8 903 1377 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=65420 $D=1
M1172 904 1374 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=51530 $D=1
M1173 905 1375 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=56160 $D=1
M1174 906 1376 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=60790 $D=1
M1175 907 1377 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=65420 $D=1
M1176 900 892 904 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=51530 $D=1
M1177 901 893 905 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=56160 $D=1
M1178 902 894 906 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=60790 $D=1
M1179 903 895 907 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=65420 $D=1
M1180 904 111 320 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=51530 $D=1
M1181 905 111 321 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=56160 $D=1
M1182 906 111 322 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=60790 $D=1
M1183 907 111 323 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=65420 $D=1
M1184 328 114 904 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=51530 $D=1
M1185 329 114 905 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=56160 $D=1
M1186 330 114 906 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=60790 $D=1
M1187 331 114 907 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=65420 $D=1
M1188 908 114 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=51530 $D=1
M1189 909 114 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=56160 $D=1
M1190 910 114 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=60790 $D=1
M1191 911 114 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=65420 $D=1
M1192 8 115 912 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=51530 $D=1
M1193 8 115 913 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=56160 $D=1
M1194 8 115 914 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=60790 $D=1
M1195 8 115 915 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=65420 $D=1
M1196 916 116 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=51530 $D=1
M1197 917 116 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=56160 $D=1
M1198 918 116 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=60790 $D=1
M1199 919 116 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=65420 $D=1
M1200 920 115 300 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=51530 $D=1
M1201 921 115 301 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=56160 $D=1
M1202 922 115 302 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=60790 $D=1
M1203 923 115 303 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=65420 $D=1
M1204 8 920 1378 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=51530 $D=1
M1205 8 921 1379 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=56160 $D=1
M1206 8 922 1380 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=60790 $D=1
M1207 8 923 1381 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=65420 $D=1
M1208 924 1378 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=51530 $D=1
M1209 925 1379 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=56160 $D=1
M1210 926 1380 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=60790 $D=1
M1211 927 1381 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=65420 $D=1
M1212 920 912 924 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=51530 $D=1
M1213 921 913 925 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=56160 $D=1
M1214 922 914 926 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=60790 $D=1
M1215 923 915 927 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=65420 $D=1
M1216 924 116 320 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=51530 $D=1
M1217 925 116 321 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=56160 $D=1
M1218 926 116 322 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=60790 $D=1
M1219 927 116 323 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=65420 $D=1
M1220 328 120 924 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=51530 $D=1
M1221 329 120 925 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=56160 $D=1
M1222 330 120 926 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=60790 $D=1
M1223 331 120 927 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=65420 $D=1
M1224 928 120 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=51530 $D=1
M1225 929 120 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=56160 $D=1
M1226 930 120 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=60790 $D=1
M1227 931 120 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=65420 $D=1
M1228 8 121 932 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=51530 $D=1
M1229 8 121 933 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=56160 $D=1
M1230 8 121 934 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=60790 $D=1
M1231 8 121 935 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=65420 $D=1
M1232 936 122 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=51530 $D=1
M1233 937 122 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=56160 $D=1
M1234 938 122 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=60790 $D=1
M1235 939 122 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=65420 $D=1
M1236 8 122 320 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=51530 $D=1
M1237 8 122 321 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=56160 $D=1
M1238 8 122 322 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=60790 $D=1
M1239 8 122 323 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=65420 $D=1
M1240 328 121 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=51530 $D=1
M1241 329 121 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=56160 $D=1
M1242 330 121 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=60790 $D=1
M1243 331 121 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=65420 $D=1
M1244 8 944 940 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=51530 $D=1
M1245 8 945 941 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=56160 $D=1
M1246 8 946 942 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=60790 $D=1
M1247 8 947 943 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=65420 $D=1
M1248 944 124 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=51530 $D=1
M1249 945 124 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=56160 $D=1
M1250 946 124 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=60790 $D=1
M1251 947 124 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=65420 $D=1
M1252 1382 320 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=51530 $D=1
M1253 1383 321 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=56160 $D=1
M1254 1384 322 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=60790 $D=1
M1255 1385 323 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=65420 $D=1
M1256 948 940 1382 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=51530 $D=1
M1257 949 941 1383 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=56160 $D=1
M1258 950 942 1384 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=60790 $D=1
M1259 951 943 1385 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=65420 $D=1
M1260 8 948 952 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=51530 $D=1
M1261 8 949 953 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=56160 $D=1
M1262 8 950 954 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=60790 $D=1
M1263 8 951 955 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=65420 $D=1
M1264 1386 952 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=51530 $D=1
M1265 1387 953 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=56160 $D=1
M1266 1388 954 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=60790 $D=1
M1267 1389 955 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=65420 $D=1
M1268 948 944 1386 8 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=51530 $D=1
M1269 949 945 1387 8 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=56160 $D=1
M1270 950 946 1388 8 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=60790 $D=1
M1271 951 947 1389 8 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=65420 $D=1
M1272 8 960 956 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=51530 $D=1
M1273 8 961 957 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=56160 $D=1
M1274 8 962 958 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=60790 $D=1
M1275 8 963 959 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=65420 $D=1
M1276 960 124 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=51530 $D=1
M1277 961 124 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=56160 $D=1
M1278 962 124 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=60790 $D=1
M1279 963 124 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=65420 $D=1
M1280 1390 328 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=51530 $D=1
M1281 1391 329 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=56160 $D=1
M1282 1392 330 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=60790 $D=1
M1283 1393 331 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=65420 $D=1
M1284 964 956 1390 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=51530 $D=1
M1285 965 957 1391 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=56160 $D=1
M1286 966 958 1392 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=60790 $D=1
M1287 967 959 1393 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=65420 $D=1
M1288 8 964 128 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=51530 $D=1
M1289 8 965 129 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=56160 $D=1
M1290 8 966 130 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=60790 $D=1
M1291 8 967 131 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=65420 $D=1
M1292 1394 128 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=51530 $D=1
M1293 1395 129 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=56160 $D=1
M1294 1396 130 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=60790 $D=1
M1295 1397 131 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=65420 $D=1
M1296 964 960 1394 8 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=51530 $D=1
M1297 965 961 1395 8 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=56160 $D=1
M1298 966 962 1396 8 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=60790 $D=1
M1299 967 963 1397 8 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=65420 $D=1
M1300 968 132 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=51530 $D=1
M1301 969 132 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=56160 $D=1
M1302 970 132 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=60790 $D=1
M1303 971 132 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=65420 $D=1
M1304 972 968 952 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=51530 $D=1
M1305 973 969 953 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=56160 $D=1
M1306 974 970 954 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=60790 $D=1
M1307 975 971 955 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=65420 $D=1
M1308 133 132 972 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=51530 $D=1
M1309 134 132 973 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=56160 $D=1
M1310 135 132 974 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=60790 $D=1
M1311 136 132 975 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=65420 $D=1
M1312 976 137 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=51530 $D=1
M1313 977 137 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=56160 $D=1
M1314 978 137 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=60790 $D=1
M1315 979 137 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=65420 $D=1
M1316 980 976 128 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=51530 $D=1
M1317 981 977 129 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=56160 $D=1
M1318 982 978 130 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=60790 $D=1
M1319 983 979 131 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=65420 $D=1
M1320 1398 137 980 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=51530 $D=1
M1321 1399 137 981 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=56160 $D=1
M1322 1400 137 982 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=60790 $D=1
M1323 1401 137 983 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=65420 $D=1
M1324 8 128 1398 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=51530 $D=1
M1325 8 129 1399 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=56160 $D=1
M1326 8 130 1400 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=60790 $D=1
M1327 8 131 1401 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=65420 $D=1
M1328 984 138 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=51530 $D=1
M1329 985 138 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=56160 $D=1
M1330 986 138 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=60790 $D=1
M1331 987 138 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=65420 $D=1
M1332 988 984 980 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=51530 $D=1
M1333 989 985 981 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=56160 $D=1
M1334 990 986 982 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=60790 $D=1
M1335 991 987 983 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=65420 $D=1
M1336 13 138 988 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=51530 $D=1
M1337 14 138 989 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=56160 $D=1
M1338 15 138 990 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=60790 $D=1
M1339 16 138 991 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=65420 $D=1
M1340 995 992 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=51530 $D=1
M1341 996 993 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=56160 $D=1
M1342 997 994 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=60790 $D=1
M1343 998 139 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=65420 $D=1
M1344 8 1003 999 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=51530 $D=1
M1345 8 1004 1000 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=56160 $D=1
M1346 8 1005 1001 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=60790 $D=1
M1347 8 1006 1002 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=65420 $D=1
M1348 1007 972 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=51530 $D=1
M1349 1008 973 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=56160 $D=1
M1350 1009 974 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=60790 $D=1
M1351 1010 975 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=65420 $D=1
M1352 1003 1007 992 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=51530 $D=1
M1353 1004 1008 993 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=56160 $D=1
M1354 1005 1009 994 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=60790 $D=1
M1355 1006 1010 139 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=65420 $D=1
M1356 995 972 1003 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=51530 $D=1
M1357 996 973 1004 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=56160 $D=1
M1358 997 974 1005 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=60790 $D=1
M1359 998 975 1006 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=65420 $D=1
M1360 1011 999 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=51530 $D=1
M1361 1012 1000 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=56160 $D=1
M1362 1013 1001 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=60790 $D=1
M1363 1014 1002 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=65420 $D=1
M1364 140 1011 988 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=51530 $D=1
M1365 992 1012 989 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=56160 $D=1
M1366 993 1013 990 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=60790 $D=1
M1367 994 1014 991 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=65420 $D=1
M1368 972 999 140 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=51530 $D=1
M1369 973 1000 992 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=56160 $D=1
M1370 974 1001 993 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=60790 $D=1
M1371 975 1002 994 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=65420 $D=1
M1372 1015 140 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=51530 $D=1
M1373 1016 992 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=56160 $D=1
M1374 1017 993 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=60790 $D=1
M1375 1018 994 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=65420 $D=1
M1376 1019 999 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=51530 $D=1
M1377 1020 1000 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=56160 $D=1
M1378 1021 1001 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=60790 $D=1
M1379 1022 1002 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=65420 $D=1
M1380 1023 1019 1015 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=51530 $D=1
M1381 1024 1020 1016 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=56160 $D=1
M1382 1025 1021 1017 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=60790 $D=1
M1383 1026 1022 1018 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=65420 $D=1
M1384 988 999 1023 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=51530 $D=1
M1385 989 1000 1024 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=56160 $D=1
M1386 990 1001 1025 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=60790 $D=1
M1387 991 1002 1026 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=65420 $D=1
M1388 1027 972 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=51530 $D=1
M1389 1028 973 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=56160 $D=1
M1390 1029 974 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=60790 $D=1
M1391 1030 975 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=65420 $D=1
M1392 8 988 1027 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=51530 $D=1
M1393 8 989 1028 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=56160 $D=1
M1394 8 990 1029 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=60790 $D=1
M1395 8 991 1030 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=65420 $D=1
M1396 1031 1023 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=51530 $D=1
M1397 1032 1024 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=56160 $D=1
M1398 1033 1025 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=60790 $D=1
M1399 1034 1026 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=65420 $D=1
M1400 1438 972 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=51530 $D=1
M1401 1439 973 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=56160 $D=1
M1402 1440 974 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=60790 $D=1
M1403 1441 975 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=65420 $D=1
M1404 1035 988 1438 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=51530 $D=1
M1405 1036 989 1439 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=56160 $D=1
M1406 1037 990 1440 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=60790 $D=1
M1407 1038 991 1441 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=65420 $D=1
M1408 1442 972 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=51530 $D=1
M1409 1443 973 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=56160 $D=1
M1410 1444 974 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=60790 $D=1
M1411 1445 975 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=65420 $D=1
M1412 1039 988 1442 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=51530 $D=1
M1413 1040 989 1443 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=56160 $D=1
M1414 1041 990 1444 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=60790 $D=1
M1415 1042 991 1445 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=65420 $D=1
M1416 1047 972 1043 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=51530 $D=1
M1417 1048 973 1044 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=56160 $D=1
M1418 1049 974 1045 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=60790 $D=1
M1419 1050 975 1046 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=65420 $D=1
M1420 1043 988 1047 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=51530 $D=1
M1421 1044 989 1048 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=56160 $D=1
M1422 1045 990 1049 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=60790 $D=1
M1423 1046 991 1050 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=65420 $D=1
M1424 8 1039 1043 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=51530 $D=1
M1425 8 1040 1044 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=56160 $D=1
M1426 8 1041 1045 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=60790 $D=1
M1427 8 1042 1046 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=65420 $D=1
M1428 1051 144 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=51530 $D=1
M1429 1052 144 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=56160 $D=1
M1430 1053 144 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=60790 $D=1
M1431 1054 144 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=65420 $D=1
M1432 1055 1051 1027 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=51530 $D=1
M1433 1056 1052 1028 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=56160 $D=1
M1434 1057 1053 1029 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=60790 $D=1
M1435 1058 1054 1030 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=65420 $D=1
M1436 1035 144 1055 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=51530 $D=1
M1437 1036 144 1056 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=56160 $D=1
M1438 1037 144 1057 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=60790 $D=1
M1439 1038 144 1058 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=65420 $D=1
M1440 1059 1051 1031 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=51530 $D=1
M1441 1060 1052 1032 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=56160 $D=1
M1442 1061 1053 1033 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=60790 $D=1
M1443 1062 1054 1034 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=65420 $D=1
M1444 1047 144 1059 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=51530 $D=1
M1445 1048 144 1060 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=56160 $D=1
M1446 1049 144 1061 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=60790 $D=1
M1447 1050 144 1062 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=65420 $D=1
M1448 1063 145 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=51530 $D=1
M1449 1064 145 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=56160 $D=1
M1450 1065 145 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=60790 $D=1
M1451 1066 145 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=65420 $D=1
M1452 1067 1063 1059 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=51530 $D=1
M1453 1068 1064 1060 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=56160 $D=1
M1454 1069 1065 1061 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=60790 $D=1
M1455 1070 1066 1062 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=65420 $D=1
M1456 1055 145 1067 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=51530 $D=1
M1457 1056 145 1068 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=56160 $D=1
M1458 1057 145 1069 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=60790 $D=1
M1459 1058 145 1070 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=65420 $D=1
M1460 17 1067 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=51530 $D=1
M1461 18 1068 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=56160 $D=1
M1462 19 1069 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=60790 $D=1
M1463 20 1070 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=65420 $D=1
M1464 1071 146 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=51530 $D=1
M1465 1072 146 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=56160 $D=1
M1466 1073 146 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=60790 $D=1
M1467 1074 146 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=65420 $D=1
M1468 1077 1071 1075 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=51530 $D=1
M1469 1078 1072 1076 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=56160 $D=1
M1470 1079 1073 147 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=60790 $D=1
M1471 1080 1074 148 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=65420 $D=1
M1472 149 146 1077 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=51530 $D=1
M1473 150 146 1078 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=56160 $D=1
M1474 1075 146 1079 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=60790 $D=1
M1475 1076 146 1080 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=65420 $D=1
M1476 1081 146 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=51530 $D=1
M1477 1082 146 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=56160 $D=1
M1478 1083 146 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=60790 $D=1
M1479 1084 146 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=65420 $D=1
M1480 1085 1081 151 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=51530 $D=1
M1481 1086 1082 152 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=56160 $D=1
M1482 1087 1083 153 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=60790 $D=1
M1483 1088 1084 154 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=65420 $D=1
M1484 155 146 1085 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=51530 $D=1
M1485 156 146 1086 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=56160 $D=1
M1486 157 146 1087 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=60790 $D=1
M1487 158 146 1088 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=65420 $D=1
M1488 1089 146 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=51530 $D=1
M1489 1090 146 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=56160 $D=1
M1490 1091 146 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=60790 $D=1
M1491 1092 146 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=65420 $D=1
M1492 1093 1089 141 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=51530 $D=1
M1493 1094 1090 143 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=56160 $D=1
M1494 1095 1091 142 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=60790 $D=1
M1495 1096 1092 159 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=65420 $D=1
M1496 160 146 1093 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=51530 $D=1
M1497 118 146 1094 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=56160 $D=1
M1498 119 146 1095 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=60790 $D=1
M1499 123 146 1096 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=65420 $D=1
M1500 1097 146 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=51530 $D=1
M1501 1098 146 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=56160 $D=1
M1502 1099 146 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=60790 $D=1
M1503 1100 146 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=65420 $D=1
M1504 1101 1097 161 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=51530 $D=1
M1505 1102 1098 162 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=56160 $D=1
M1506 1103 1099 163 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=60790 $D=1
M1507 1104 1100 164 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=65420 $D=1
M1508 165 146 1101 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=51530 $D=1
M1509 166 146 1102 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=56160 $D=1
M1510 167 146 1103 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=60790 $D=1
M1511 168 146 1104 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=65420 $D=1
M1512 1105 146 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=51530 $D=1
M1513 1106 146 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=56160 $D=1
M1514 1107 146 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=60790 $D=1
M1515 1108 146 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=65420 $D=1
M1516 1109 1105 169 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=51530 $D=1
M1517 1110 1106 170 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=56160 $D=1
M1518 1111 1107 171 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=60790 $D=1
M1519 1112 1108 172 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=65420 $D=1
M1520 173 146 1109 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=51530 $D=1
M1521 173 146 1110 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=56160 $D=1
M1522 173 146 1111 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=60790 $D=1
M1523 173 146 1112 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=65420 $D=1
M1524 8 972 1402 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=51530 $D=1
M1525 8 973 1403 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=56160 $D=1
M1526 8 974 1404 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=60790 $D=1
M1527 8 975 1405 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=65420 $D=1
M1528 150 1402 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=51530 $D=1
M1529 1075 1403 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=56160 $D=1
M1530 1076 1404 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=60790 $D=1
M1531 147 1405 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=65420 $D=1
M1532 1113 174 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=51530 $D=1
M1533 1114 174 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=56160 $D=1
M1534 1115 174 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=60790 $D=1
M1535 1116 174 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=65420 $D=1
M1536 157 1113 150 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=51530 $D=1
M1537 158 1114 1075 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=56160 $D=1
M1538 151 1115 1076 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=60790 $D=1
M1539 152 1116 147 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=65420 $D=1
M1540 1077 174 157 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=51530 $D=1
M1541 1078 174 158 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=56160 $D=1
M1542 1079 174 151 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=60790 $D=1
M1543 1080 174 152 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=65420 $D=1
M1544 1117 175 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=51530 $D=1
M1545 1118 175 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=56160 $D=1
M1546 1119 175 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=60790 $D=1
M1547 1120 175 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=65420 $D=1
M1548 176 1117 157 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=51530 $D=1
M1549 125 1118 158 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=56160 $D=1
M1550 126 1119 151 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=60790 $D=1
M1551 127 1120 152 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=65420 $D=1
M1552 1085 175 176 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=51530 $D=1
M1553 1086 175 125 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=56160 $D=1
M1554 1087 175 126 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=60790 $D=1
M1555 1088 175 127 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=65420 $D=1
M1556 1121 177 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=51530 $D=1
M1557 1122 177 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=56160 $D=1
M1558 1123 177 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=60790 $D=1
M1559 1124 177 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=65420 $D=1
M1560 178 1121 176 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=51530 $D=1
M1561 112 1122 125 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=56160 $D=1
M1562 113 1123 126 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=60790 $D=1
M1563 117 1124 127 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=65420 $D=1
M1564 1093 177 178 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=51530 $D=1
M1565 1094 177 112 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=56160 $D=1
M1566 1095 177 113 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=60790 $D=1
M1567 1096 177 117 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=65420 $D=1
M1568 1125 179 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=51530 $D=1
M1569 1126 179 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=56160 $D=1
M1570 1127 179 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=60790 $D=1
M1571 1128 179 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=65420 $D=1
M1572 180 1125 178 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=51530 $D=1
M1573 181 1126 112 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=56160 $D=1
M1574 182 1127 113 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=60790 $D=1
M1575 183 1128 117 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=65420 $D=1
M1576 1101 179 180 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=51530 $D=1
M1577 1102 179 181 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=56160 $D=1
M1578 1103 179 182 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=60790 $D=1
M1579 1104 179 183 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=65420 $D=1
M1580 1129 184 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=51530 $D=1
M1581 1130 184 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=56160 $D=1
M1582 1131 184 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=60790 $D=1
M1583 1132 184 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=65420 $D=1
M1584 272 1129 180 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=51530 $D=1
M1585 273 1130 181 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=56160 $D=1
M1586 274 1131 182 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=60790 $D=1
M1587 275 1132 183 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=65420 $D=1
M1588 1109 184 272 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=51530 $D=1
M1589 1110 184 273 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=56160 $D=1
M1590 1111 184 274 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=60790 $D=1
M1591 1112 184 275 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=65420 $D=1
M1592 1133 185 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=51530 $D=1
M1593 1134 185 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=56160 $D=1
M1594 1135 185 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=60790 $D=1
M1595 1136 185 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=65420 $D=1
M1596 1137 1133 128 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=51530 $D=1
M1597 1138 1134 129 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=56160 $D=1
M1598 1139 1135 130 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=60790 $D=1
M1599 1140 1136 131 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=65420 $D=1
M1600 13 185 1137 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=51530 $D=1
M1601 14 185 1138 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=56160 $D=1
M1602 15 185 1139 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=60790 $D=1
M1603 16 185 1140 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=65420 $D=1
M1604 1446 952 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=51530 $D=1
M1605 1447 953 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=56160 $D=1
M1606 1448 954 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=60790 $D=1
M1607 1449 955 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=65420 $D=1
M1608 1141 1137 1446 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=51530 $D=1
M1609 1142 1138 1447 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=56160 $D=1
M1610 1143 1139 1448 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=60790 $D=1
M1611 1144 1140 1449 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=65420 $D=1
M1612 1149 952 1145 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=51530 $D=1
M1613 1150 953 1146 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=56160 $D=1
M1614 1151 954 1147 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=60790 $D=1
M1615 1152 955 1148 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=65420 $D=1
M1616 1145 1137 1149 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=51530 $D=1
M1617 1146 1138 1150 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=56160 $D=1
M1618 1147 1139 1151 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=60790 $D=1
M1619 1148 1140 1152 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=65420 $D=1
M1620 8 1141 1145 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=51530 $D=1
M1621 8 1142 1146 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=56160 $D=1
M1622 8 1143 1147 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=60790 $D=1
M1623 8 1144 1148 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=65420 $D=1
M1624 1450 186 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=51530 $D=1
M1625 1451 1153 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=56160 $D=1
M1626 1452 1154 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=60790 $D=1
M1627 1453 1155 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=65420 $D=1
M1628 1406 1149 1450 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=51530 $D=1
M1629 1407 1150 1451 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=56160 $D=1
M1630 1408 1151 1452 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=60790 $D=1
M1631 1409 1152 1453 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=65420 $D=1
M1632 1153 1406 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=51530 $D=1
M1633 1154 1407 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=56160 $D=1
M1634 1155 1408 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=60790 $D=1
M1635 187 1409 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=65420 $D=1
M1636 1156 952 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=51530 $D=1
M1637 1157 953 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=56160 $D=1
M1638 1158 954 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=60790 $D=1
M1639 1159 955 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=65420 $D=1
M1640 8 1160 1156 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=51530 $D=1
M1641 8 1161 1157 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=56160 $D=1
M1642 8 1162 1158 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=60790 $D=1
M1643 8 1163 1159 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=65420 $D=1
M1644 1160 1137 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=51530 $D=1
M1645 1161 1138 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=56160 $D=1
M1646 1162 1139 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=60790 $D=1
M1647 1163 1140 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=65420 $D=1
M1648 1454 1156 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=51530 $D=1
M1649 1455 1157 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=56160 $D=1
M1650 1456 1158 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=60790 $D=1
M1651 1457 1159 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=65420 $D=1
M1652 1164 186 1454 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=51530 $D=1
M1653 1165 1153 1455 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=56160 $D=1
M1654 1166 1154 1456 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=60790 $D=1
M1655 1167 1155 1457 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=65420 $D=1
M1656 1171 188 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=51530 $D=1
M1657 1172 1168 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=56160 $D=1
M1658 1173 1169 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=60790 $D=1
M1659 1174 1170 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=65420 $D=1
M1660 1458 1164 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=51530 $D=1
M1661 1459 1165 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=56160 $D=1
M1662 1460 1166 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=60790 $D=1
M1663 1461 1167 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=65420 $D=1
M1664 1168 1171 1458 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=51530 $D=1
M1665 1169 1172 1459 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=56160 $D=1
M1666 1170 1173 1460 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=60790 $D=1
M1667 189 1174 1461 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=65420 $D=1
M1668 1178 1175 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=51530 $D=1
M1669 1179 1176 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=56160 $D=1
M1670 1180 1177 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=60790 $D=1
M1671 1181 190 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=65420 $D=1
M1672 8 1186 1182 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=51530 $D=1
M1673 8 1187 1183 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=56160 $D=1
M1674 8 1188 1184 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=60790 $D=1
M1675 8 1189 1185 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=65420 $D=1
M1676 1190 133 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=51530 $D=1
M1677 1191 134 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=56160 $D=1
M1678 1192 135 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=60790 $D=1
M1679 1193 136 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=65420 $D=1
M1680 1186 1190 1175 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=51530 $D=1
M1681 1187 1191 1176 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=56160 $D=1
M1682 1188 1192 1177 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=60790 $D=1
M1683 1189 1193 190 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=65420 $D=1
M1684 1178 133 1186 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=51530 $D=1
M1685 1179 134 1187 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=56160 $D=1
M1686 1180 135 1188 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=60790 $D=1
M1687 1181 136 1189 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=65420 $D=1
M1688 1194 1182 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=51530 $D=1
M1689 1195 1183 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=56160 $D=1
M1690 1196 1184 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=60790 $D=1
M1691 1197 1185 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=65420 $D=1
M1692 191 1194 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=51530 $D=1
M1693 1175 1195 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=56160 $D=1
M1694 1176 1196 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=60790 $D=1
M1695 1177 1197 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=65420 $D=1
M1696 133 1182 191 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=51530 $D=1
M1697 134 1183 1175 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=56160 $D=1
M1698 135 1184 1176 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=60790 $D=1
M1699 136 1185 1177 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=65420 $D=1
M1700 1198 191 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=51530 $D=1
M1701 1199 1175 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=56160 $D=1
M1702 1200 1176 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=60790 $D=1
M1703 1201 1177 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=65420 $D=1
M1704 1202 1182 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=51530 $D=1
M1705 1203 1183 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=56160 $D=1
M1706 1204 1184 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=60790 $D=1
M1707 1205 1185 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=65420 $D=1
M1708 276 1202 1198 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=51530 $D=1
M1709 277 1203 1199 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=56160 $D=1
M1710 278 1204 1200 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=60790 $D=1
M1711 279 1205 1201 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=65420 $D=1
M1712 8 1182 276 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=51530 $D=1
M1713 8 1183 277 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=56160 $D=1
M1714 8 1184 278 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=60790 $D=1
M1715 8 1185 279 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=65420 $D=1
M1716 1206 192 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=51530 $D=1
M1717 1207 192 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=56160 $D=1
M1718 1208 192 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=60790 $D=1
M1719 1209 192 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=65420 $D=1
M1720 1210 1206 276 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=51530 $D=1
M1721 1211 1207 277 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=56160 $D=1
M1722 1212 1208 278 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=60790 $D=1
M1723 1213 1209 279 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=65420 $D=1
M1724 17 192 1210 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=51530 $D=1
M1725 18 192 1211 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=56160 $D=1
M1726 19 192 1212 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=60790 $D=1
M1727 20 192 1213 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=65420 $D=1
M1728 1214 193 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=51530 $D=1
M1729 1215 193 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=56160 $D=1
M1730 1216 193 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=60790 $D=1
M1731 1217 193 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=65420 $D=1
M1732 1218 1214 1210 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=51530 $D=1
M1733 1219 1215 1211 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=56160 $D=1
M1734 1220 1216 1212 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=60790 $D=1
M1735 1221 1217 1213 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=65420 $D=1
M1736 8 193 1218 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=51530 $D=1
M1737 8 193 1219 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=56160 $D=1
M1738 8 193 1220 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=60790 $D=1
M1739 8 193 1221 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=65420 $D=1
M1740 1222 124 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=51530 $D=1
M1741 1223 124 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=56160 $D=1
M1742 1224 124 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=60790 $D=1
M1743 1225 124 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=65420 $D=1
M1744 8 1222 1226 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=51530 $D=1
M1745 8 1223 1227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=56160 $D=1
M1746 8 1224 1228 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=60790 $D=1
M1747 8 1225 1229 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=65420 $D=1
M1748 1230 124 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=51530 $D=1
M1749 1231 124 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=56160 $D=1
M1750 1232 124 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=60790 $D=1
M1751 1233 124 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=65420 $D=1
M1752 1234 1222 1218 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=51530 $D=1
M1753 1235 1223 1219 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=56160 $D=1
M1754 1236 1224 1220 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=60790 $D=1
M1755 1237 1225 1221 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=65420 $D=1
M1756 8 1234 1410 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=51530 $D=1
M1757 8 1235 1411 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=56160 $D=1
M1758 8 1236 1412 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=60790 $D=1
M1759 8 1237 1413 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=65420 $D=1
M1760 1238 1410 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=51530 $D=1
M1761 1239 1411 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=56160 $D=1
M1762 1240 1412 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=60790 $D=1
M1763 1241 1413 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=65420 $D=1
M1764 1234 1226 1238 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=51530 $D=1
M1765 1235 1227 1239 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=56160 $D=1
M1766 1236 1228 1240 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=60790 $D=1
M1767 1237 1229 1241 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=65420 $D=1
M1768 1242 124 1238 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=51530 $D=1
M1769 1243 124 1239 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=56160 $D=1
M1770 1244 124 1240 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=60790 $D=1
M1771 1245 124 1241 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=65420 $D=1
M1772 8 1250 1246 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=51530 $D=1
M1773 8 1251 1247 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=56160 $D=1
M1774 8 1252 1248 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=60790 $D=1
M1775 8 1253 1249 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=65420 $D=1
M1776 1250 124 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=51530 $D=1
M1777 1251 124 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=56160 $D=1
M1778 1252 124 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=60790 $D=1
M1779 1253 124 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=65420 $D=1
M1780 1414 1242 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=51530 $D=1
M1781 1415 1243 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=56160 $D=1
M1782 1416 1244 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=60790 $D=1
M1783 1417 1245 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=65420 $D=1
M1784 1254 1246 1414 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=51530 $D=1
M1785 1255 1247 1415 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=56160 $D=1
M1786 1256 1248 1416 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=60790 $D=1
M1787 1257 1249 1417 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=65420 $D=1
M1788 8 1254 133 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=51530 $D=1
M1789 8 1255 134 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=56160 $D=1
M1790 8 1256 135 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=60790 $D=1
M1791 8 1257 136 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=65420 $D=1
M1792 1418 133 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=51530 $D=1
M1793 1419 134 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=56160 $D=1
M1794 1420 135 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=60790 $D=1
M1795 1421 136 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=65420 $D=1
M1796 1254 1250 1418 8 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=51530 $D=1
M1797 1255 1251 1419 8 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=56160 $D=1
M1798 1256 1252 1420 8 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=60790 $D=1
M1799 1257 1253 1421 8 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=65420 $D=1
M1800 224 1 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=52780 $D=0
M1801 225 1 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=57410 $D=0
M1802 226 1 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=62040 $D=0
M1803 227 1 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=66670 $D=0
M1804 228 1 2 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=52780 $D=0
M1805 229 1 3 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=57410 $D=0
M1806 230 1 4 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=62040 $D=0
M1807 231 1 5 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=66670 $D=0
M1808 8 224 228 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=52780 $D=0
M1809 8 225 229 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=57410 $D=0
M1810 8 226 230 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=62040 $D=0
M1811 8 227 231 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=66670 $D=0
M1812 232 1 6 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=52780 $D=0
M1813 233 1 6 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=57410 $D=0
M1814 234 1 6 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=62040 $D=0
M1815 235 1 6 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=66670 $D=0
M1816 7 224 232 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=52780 $D=0
M1817 7 225 233 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=57410 $D=0
M1818 7 226 234 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=62040 $D=0
M1819 7 227 235 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=66670 $D=0
M1820 236 1 8 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=52780 $D=0
M1821 237 1 8 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=57410 $D=0
M1822 238 1 8 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=62040 $D=0
M1823 239 1 8 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=66670 $D=0
M1824 8 224 236 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=52780 $D=0
M1825 8 225 237 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=57410 $D=0
M1826 8 226 238 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=62040 $D=0
M1827 8 227 239 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=66670 $D=0
M1828 244 9 236 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=52780 $D=0
M1829 245 9 237 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=57410 $D=0
M1830 246 9 238 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=62040 $D=0
M1831 247 9 239 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=66670 $D=0
M1832 240 9 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=52780 $D=0
M1833 241 9 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=57410 $D=0
M1834 242 9 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=62040 $D=0
M1835 243 9 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=66670 $D=0
M1836 248 9 232 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=52780 $D=0
M1837 249 9 233 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=57410 $D=0
M1838 250 9 234 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=62040 $D=0
M1839 251 9 235 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=66670 $D=0
M1840 228 240 248 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=52780 $D=0
M1841 229 241 249 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=57410 $D=0
M1842 230 242 250 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=62040 $D=0
M1843 231 243 251 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=66670 $D=0
M1844 252 10 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=52780 $D=0
M1845 253 10 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=57410 $D=0
M1846 254 10 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=62040 $D=0
M1847 255 10 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=66670 $D=0
M1848 256 10 248 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=52780 $D=0
M1849 257 10 249 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=57410 $D=0
M1850 258 10 250 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=62040 $D=0
M1851 259 10 251 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=66670 $D=0
M1852 244 252 256 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=52780 $D=0
M1853 245 253 257 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=57410 $D=0
M1854 246 254 258 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=62040 $D=0
M1855 247 255 259 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=66670 $D=0
M1856 260 12 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=52780 $D=0
M1857 261 12 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=57410 $D=0
M1858 262 12 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=62040 $D=0
M1859 263 12 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=66670 $D=0
M1860 264 12 8 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=52780 $D=0
M1861 265 12 8 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=57410 $D=0
M1862 266 12 8 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=62040 $D=0
M1863 267 12 8 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=66670 $D=0
M1864 13 260 264 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=52780 $D=0
M1865 14 261 265 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=57410 $D=0
M1866 15 262 266 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=62040 $D=0
M1867 16 263 267 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=66670 $D=0
M1868 268 12 17 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=52780 $D=0
M1869 269 12 18 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=57410 $D=0
M1870 270 12 19 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=62040 $D=0
M1871 271 12 20 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=66670 $D=0
M1872 272 260 268 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=52780 $D=0
M1873 273 261 269 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=57410 $D=0
M1874 274 262 270 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=62040 $D=0
M1875 275 263 271 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=66670 $D=0
M1876 280 12 276 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=52780 $D=0
M1877 281 12 277 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=57410 $D=0
M1878 282 12 278 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=62040 $D=0
M1879 283 12 279 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=66670 $D=0
M1880 256 260 280 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=52780 $D=0
M1881 257 261 281 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=57410 $D=0
M1882 258 262 282 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=62040 $D=0
M1883 259 263 283 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=66670 $D=0
M1884 288 21 280 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=52780 $D=0
M1885 289 21 281 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=57410 $D=0
M1886 290 21 282 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=62040 $D=0
M1887 291 21 283 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=66670 $D=0
M1888 284 21 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=52780 $D=0
M1889 285 21 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=57410 $D=0
M1890 286 21 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=62040 $D=0
M1891 287 21 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=66670 $D=0
M1892 292 21 268 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=52780 $D=0
M1893 293 21 269 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=57410 $D=0
M1894 294 21 270 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=62040 $D=0
M1895 295 21 271 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=66670 $D=0
M1896 264 284 292 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=52780 $D=0
M1897 265 285 293 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=57410 $D=0
M1898 266 286 294 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=62040 $D=0
M1899 267 287 295 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=66670 $D=0
M1900 296 22 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=52780 $D=0
M1901 297 22 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=57410 $D=0
M1902 298 22 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=62040 $D=0
M1903 299 22 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=66670 $D=0
M1904 300 22 292 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=52780 $D=0
M1905 301 22 293 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=57410 $D=0
M1906 302 22 294 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=62040 $D=0
M1907 303 22 295 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=66670 $D=0
M1908 288 296 300 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=52780 $D=0
M1909 289 297 301 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=57410 $D=0
M1910 290 298 302 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=62040 $D=0
M1911 291 299 303 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=66670 $D=0
M1912 11 23 304 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=52780 $D=0
M1913 11 23 305 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=57410 $D=0
M1914 11 23 306 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=62040 $D=0
M1915 11 23 307 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=66670 $D=0
M1916 308 24 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=52780 $D=0
M1917 309 24 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=57410 $D=0
M1918 310 24 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=62040 $D=0
M1919 311 24 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=66670 $D=0
M1920 312 304 300 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=52780 $D=0
M1921 313 305 301 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=57410 $D=0
M1922 314 306 302 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=62040 $D=0
M1923 315 307 303 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=66670 $D=0
M1924 11 312 1258 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=52780 $D=0
M1925 11 313 1259 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=57410 $D=0
M1926 11 314 1260 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=62040 $D=0
M1927 11 315 1261 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=66670 $D=0
M1928 316 1258 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=52780 $D=0
M1929 317 1259 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=57410 $D=0
M1930 318 1260 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=62040 $D=0
M1931 319 1261 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=66670 $D=0
M1932 312 23 316 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=52780 $D=0
M1933 313 23 317 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=57410 $D=0
M1934 314 23 318 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=62040 $D=0
M1935 315 23 319 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=66670 $D=0
M1936 316 308 320 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=52780 $D=0
M1937 317 309 321 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=57410 $D=0
M1938 318 310 322 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=62040 $D=0
M1939 319 311 323 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=66670 $D=0
M1940 328 324 316 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=52780 $D=0
M1941 329 325 317 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=57410 $D=0
M1942 330 326 318 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=62040 $D=0
M1943 331 327 319 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=66670 $D=0
M1944 324 25 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=52780 $D=0
M1945 325 25 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=57410 $D=0
M1946 326 25 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=62040 $D=0
M1947 327 25 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=66670 $D=0
M1948 11 26 332 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=52780 $D=0
M1949 11 26 333 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=57410 $D=0
M1950 11 26 334 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=62040 $D=0
M1951 11 26 335 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=66670 $D=0
M1952 336 27 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=52780 $D=0
M1953 337 27 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=57410 $D=0
M1954 338 27 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=62040 $D=0
M1955 339 27 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=66670 $D=0
M1956 340 332 300 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=52780 $D=0
M1957 341 333 301 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=57410 $D=0
M1958 342 334 302 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=62040 $D=0
M1959 343 335 303 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=66670 $D=0
M1960 11 340 1262 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=52780 $D=0
M1961 11 341 1263 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=57410 $D=0
M1962 11 342 1264 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=62040 $D=0
M1963 11 343 1265 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=66670 $D=0
M1964 344 1262 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=52780 $D=0
M1965 345 1263 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=57410 $D=0
M1966 346 1264 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=62040 $D=0
M1967 347 1265 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=66670 $D=0
M1968 340 26 344 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=52780 $D=0
M1969 341 26 345 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=57410 $D=0
M1970 342 26 346 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=62040 $D=0
M1971 343 26 347 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=66670 $D=0
M1972 344 336 320 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=52780 $D=0
M1973 345 337 321 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=57410 $D=0
M1974 346 338 322 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=62040 $D=0
M1975 347 339 323 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=66670 $D=0
M1976 328 348 344 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=52780 $D=0
M1977 329 349 345 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=57410 $D=0
M1978 330 350 346 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=62040 $D=0
M1979 331 351 347 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=66670 $D=0
M1980 348 28 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=52780 $D=0
M1981 349 28 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=57410 $D=0
M1982 350 28 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=62040 $D=0
M1983 351 28 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=66670 $D=0
M1984 11 29 352 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=52780 $D=0
M1985 11 29 353 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=57410 $D=0
M1986 11 29 354 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=62040 $D=0
M1987 11 29 355 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=66670 $D=0
M1988 356 30 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=52780 $D=0
M1989 357 30 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=57410 $D=0
M1990 358 30 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=62040 $D=0
M1991 359 30 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=66670 $D=0
M1992 360 352 300 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=52780 $D=0
M1993 361 353 301 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=57410 $D=0
M1994 362 354 302 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=62040 $D=0
M1995 363 355 303 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=66670 $D=0
M1996 11 360 1266 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=52780 $D=0
M1997 11 361 1267 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=57410 $D=0
M1998 11 362 1268 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=62040 $D=0
M1999 11 363 1269 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=66670 $D=0
M2000 364 1266 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=52780 $D=0
M2001 365 1267 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=57410 $D=0
M2002 366 1268 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=62040 $D=0
M2003 367 1269 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=66670 $D=0
M2004 360 29 364 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=52780 $D=0
M2005 361 29 365 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=57410 $D=0
M2006 362 29 366 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=62040 $D=0
M2007 363 29 367 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=66670 $D=0
M2008 364 356 320 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=52780 $D=0
M2009 365 357 321 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=57410 $D=0
M2010 366 358 322 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=62040 $D=0
M2011 367 359 323 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=66670 $D=0
M2012 328 368 364 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=52780 $D=0
M2013 329 369 365 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=57410 $D=0
M2014 330 370 366 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=62040 $D=0
M2015 331 371 367 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=66670 $D=0
M2016 368 31 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=52780 $D=0
M2017 369 31 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=57410 $D=0
M2018 370 31 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=62040 $D=0
M2019 371 31 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=66670 $D=0
M2020 11 32 372 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=52780 $D=0
M2021 11 32 373 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=57410 $D=0
M2022 11 32 374 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=62040 $D=0
M2023 11 32 375 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=66670 $D=0
M2024 376 33 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=52780 $D=0
M2025 377 33 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=57410 $D=0
M2026 378 33 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=62040 $D=0
M2027 379 33 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=66670 $D=0
M2028 380 372 300 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=52780 $D=0
M2029 381 373 301 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=57410 $D=0
M2030 382 374 302 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=62040 $D=0
M2031 383 375 303 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=66670 $D=0
M2032 11 380 1270 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=52780 $D=0
M2033 11 381 1271 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=57410 $D=0
M2034 11 382 1272 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=62040 $D=0
M2035 11 383 1273 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=66670 $D=0
M2036 384 1270 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=52780 $D=0
M2037 385 1271 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=57410 $D=0
M2038 386 1272 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=62040 $D=0
M2039 387 1273 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=66670 $D=0
M2040 380 32 384 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=52780 $D=0
M2041 381 32 385 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=57410 $D=0
M2042 382 32 386 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=62040 $D=0
M2043 383 32 387 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=66670 $D=0
M2044 384 376 320 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=52780 $D=0
M2045 385 377 321 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=57410 $D=0
M2046 386 378 322 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=62040 $D=0
M2047 387 379 323 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=66670 $D=0
M2048 328 388 384 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=52780 $D=0
M2049 329 389 385 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=57410 $D=0
M2050 330 390 386 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=62040 $D=0
M2051 331 391 387 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=66670 $D=0
M2052 388 34 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=52780 $D=0
M2053 389 34 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=57410 $D=0
M2054 390 34 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=62040 $D=0
M2055 391 34 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=66670 $D=0
M2056 11 35 392 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=52780 $D=0
M2057 11 35 393 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=57410 $D=0
M2058 11 35 394 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=62040 $D=0
M2059 11 35 395 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=66670 $D=0
M2060 396 36 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=52780 $D=0
M2061 397 36 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=57410 $D=0
M2062 398 36 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=62040 $D=0
M2063 399 36 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=66670 $D=0
M2064 400 392 300 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=52780 $D=0
M2065 401 393 301 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=57410 $D=0
M2066 402 394 302 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=62040 $D=0
M2067 403 395 303 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=66670 $D=0
M2068 11 400 1274 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=52780 $D=0
M2069 11 401 1275 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=57410 $D=0
M2070 11 402 1276 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=62040 $D=0
M2071 11 403 1277 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=66670 $D=0
M2072 404 1274 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=52780 $D=0
M2073 405 1275 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=57410 $D=0
M2074 406 1276 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=62040 $D=0
M2075 407 1277 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=66670 $D=0
M2076 400 35 404 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=52780 $D=0
M2077 401 35 405 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=57410 $D=0
M2078 402 35 406 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=62040 $D=0
M2079 403 35 407 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=66670 $D=0
M2080 404 396 320 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=52780 $D=0
M2081 405 397 321 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=57410 $D=0
M2082 406 398 322 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=62040 $D=0
M2083 407 399 323 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=66670 $D=0
M2084 328 408 404 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=52780 $D=0
M2085 329 409 405 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=57410 $D=0
M2086 330 410 406 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=62040 $D=0
M2087 331 411 407 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=66670 $D=0
M2088 408 37 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=52780 $D=0
M2089 409 37 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=57410 $D=0
M2090 410 37 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=62040 $D=0
M2091 411 37 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=66670 $D=0
M2092 11 38 412 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=52780 $D=0
M2093 11 38 413 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=57410 $D=0
M2094 11 38 414 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=62040 $D=0
M2095 11 38 415 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=66670 $D=0
M2096 416 39 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=52780 $D=0
M2097 417 39 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=57410 $D=0
M2098 418 39 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=62040 $D=0
M2099 419 39 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=66670 $D=0
M2100 420 412 300 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=52780 $D=0
M2101 421 413 301 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=57410 $D=0
M2102 422 414 302 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=62040 $D=0
M2103 423 415 303 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=66670 $D=0
M2104 11 420 1278 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=52780 $D=0
M2105 11 421 1279 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=57410 $D=0
M2106 11 422 1280 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=62040 $D=0
M2107 11 423 1281 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=66670 $D=0
M2108 424 1278 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=52780 $D=0
M2109 425 1279 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=57410 $D=0
M2110 426 1280 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=62040 $D=0
M2111 427 1281 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=66670 $D=0
M2112 420 38 424 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=52780 $D=0
M2113 421 38 425 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=57410 $D=0
M2114 422 38 426 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=62040 $D=0
M2115 423 38 427 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=66670 $D=0
M2116 424 416 320 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=52780 $D=0
M2117 425 417 321 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=57410 $D=0
M2118 426 418 322 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=62040 $D=0
M2119 427 419 323 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=66670 $D=0
M2120 328 428 424 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=52780 $D=0
M2121 329 429 425 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=57410 $D=0
M2122 330 430 426 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=62040 $D=0
M2123 331 431 427 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=66670 $D=0
M2124 428 40 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=52780 $D=0
M2125 429 40 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=57410 $D=0
M2126 430 40 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=62040 $D=0
M2127 431 40 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=66670 $D=0
M2128 11 41 432 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=52780 $D=0
M2129 11 41 433 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=57410 $D=0
M2130 11 41 434 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=62040 $D=0
M2131 11 41 435 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=66670 $D=0
M2132 436 42 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=52780 $D=0
M2133 437 42 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=57410 $D=0
M2134 438 42 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=62040 $D=0
M2135 439 42 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=66670 $D=0
M2136 440 432 300 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=52780 $D=0
M2137 441 433 301 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=57410 $D=0
M2138 442 434 302 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=62040 $D=0
M2139 443 435 303 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=66670 $D=0
M2140 11 440 1282 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=52780 $D=0
M2141 11 441 1283 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=57410 $D=0
M2142 11 442 1284 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=62040 $D=0
M2143 11 443 1285 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=66670 $D=0
M2144 444 1282 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=52780 $D=0
M2145 445 1283 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=57410 $D=0
M2146 446 1284 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=62040 $D=0
M2147 447 1285 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=66670 $D=0
M2148 440 41 444 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=52780 $D=0
M2149 441 41 445 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=57410 $D=0
M2150 442 41 446 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=62040 $D=0
M2151 443 41 447 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=66670 $D=0
M2152 444 436 320 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=52780 $D=0
M2153 445 437 321 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=57410 $D=0
M2154 446 438 322 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=62040 $D=0
M2155 447 439 323 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=66670 $D=0
M2156 328 448 444 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=52780 $D=0
M2157 329 449 445 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=57410 $D=0
M2158 330 450 446 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=62040 $D=0
M2159 331 451 447 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=66670 $D=0
M2160 448 43 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=52780 $D=0
M2161 449 43 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=57410 $D=0
M2162 450 43 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=62040 $D=0
M2163 451 43 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=66670 $D=0
M2164 11 44 452 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=52780 $D=0
M2165 11 44 453 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=57410 $D=0
M2166 11 44 454 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=62040 $D=0
M2167 11 44 455 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=66670 $D=0
M2168 456 45 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=52780 $D=0
M2169 457 45 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=57410 $D=0
M2170 458 45 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=62040 $D=0
M2171 459 45 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=66670 $D=0
M2172 460 452 300 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=52780 $D=0
M2173 461 453 301 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=57410 $D=0
M2174 462 454 302 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=62040 $D=0
M2175 463 455 303 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=66670 $D=0
M2176 11 460 1286 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=52780 $D=0
M2177 11 461 1287 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=57410 $D=0
M2178 11 462 1288 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=62040 $D=0
M2179 11 463 1289 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=66670 $D=0
M2180 464 1286 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=52780 $D=0
M2181 465 1287 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=57410 $D=0
M2182 466 1288 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=62040 $D=0
M2183 467 1289 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=66670 $D=0
M2184 460 44 464 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=52780 $D=0
M2185 461 44 465 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=57410 $D=0
M2186 462 44 466 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=62040 $D=0
M2187 463 44 467 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=66670 $D=0
M2188 464 456 320 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=52780 $D=0
M2189 465 457 321 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=57410 $D=0
M2190 466 458 322 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=62040 $D=0
M2191 467 459 323 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=66670 $D=0
M2192 328 468 464 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=52780 $D=0
M2193 329 469 465 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=57410 $D=0
M2194 330 470 466 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=62040 $D=0
M2195 331 471 467 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=66670 $D=0
M2196 468 46 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=52780 $D=0
M2197 469 46 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=57410 $D=0
M2198 470 46 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=62040 $D=0
M2199 471 46 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=66670 $D=0
M2200 11 47 472 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=52780 $D=0
M2201 11 47 473 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=57410 $D=0
M2202 11 47 474 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=62040 $D=0
M2203 11 47 475 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=66670 $D=0
M2204 476 48 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=52780 $D=0
M2205 477 48 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=57410 $D=0
M2206 478 48 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=62040 $D=0
M2207 479 48 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=66670 $D=0
M2208 480 472 300 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=52780 $D=0
M2209 481 473 301 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=57410 $D=0
M2210 482 474 302 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=62040 $D=0
M2211 483 475 303 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=66670 $D=0
M2212 11 480 1290 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=52780 $D=0
M2213 11 481 1291 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=57410 $D=0
M2214 11 482 1292 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=62040 $D=0
M2215 11 483 1293 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=66670 $D=0
M2216 484 1290 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=52780 $D=0
M2217 485 1291 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=57410 $D=0
M2218 486 1292 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=62040 $D=0
M2219 487 1293 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=66670 $D=0
M2220 480 47 484 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=52780 $D=0
M2221 481 47 485 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=57410 $D=0
M2222 482 47 486 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=62040 $D=0
M2223 483 47 487 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=66670 $D=0
M2224 484 476 320 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=52780 $D=0
M2225 485 477 321 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=57410 $D=0
M2226 486 478 322 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=62040 $D=0
M2227 487 479 323 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=66670 $D=0
M2228 328 488 484 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=52780 $D=0
M2229 329 489 485 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=57410 $D=0
M2230 330 490 486 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=62040 $D=0
M2231 331 491 487 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=66670 $D=0
M2232 488 49 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=52780 $D=0
M2233 489 49 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=57410 $D=0
M2234 490 49 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=62040 $D=0
M2235 491 49 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=66670 $D=0
M2236 11 50 492 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=52780 $D=0
M2237 11 50 493 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=57410 $D=0
M2238 11 50 494 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=62040 $D=0
M2239 11 50 495 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=66670 $D=0
M2240 496 51 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=52780 $D=0
M2241 497 51 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=57410 $D=0
M2242 498 51 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=62040 $D=0
M2243 499 51 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=66670 $D=0
M2244 500 492 300 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=52780 $D=0
M2245 501 493 301 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=57410 $D=0
M2246 502 494 302 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=62040 $D=0
M2247 503 495 303 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=66670 $D=0
M2248 11 500 1294 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=52780 $D=0
M2249 11 501 1295 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=57410 $D=0
M2250 11 502 1296 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=62040 $D=0
M2251 11 503 1297 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=66670 $D=0
M2252 504 1294 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=52780 $D=0
M2253 505 1295 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=57410 $D=0
M2254 506 1296 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=62040 $D=0
M2255 507 1297 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=66670 $D=0
M2256 500 50 504 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=52780 $D=0
M2257 501 50 505 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=57410 $D=0
M2258 502 50 506 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=62040 $D=0
M2259 503 50 507 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=66670 $D=0
M2260 504 496 320 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=52780 $D=0
M2261 505 497 321 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=57410 $D=0
M2262 506 498 322 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=62040 $D=0
M2263 507 499 323 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=66670 $D=0
M2264 328 508 504 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=52780 $D=0
M2265 329 509 505 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=57410 $D=0
M2266 330 510 506 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=62040 $D=0
M2267 331 511 507 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=66670 $D=0
M2268 508 52 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=52780 $D=0
M2269 509 52 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=57410 $D=0
M2270 510 52 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=62040 $D=0
M2271 511 52 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=66670 $D=0
M2272 11 53 512 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=52780 $D=0
M2273 11 53 513 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=57410 $D=0
M2274 11 53 514 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=62040 $D=0
M2275 11 53 515 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=66670 $D=0
M2276 516 54 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=52780 $D=0
M2277 517 54 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=57410 $D=0
M2278 518 54 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=62040 $D=0
M2279 519 54 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=66670 $D=0
M2280 520 512 300 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=52780 $D=0
M2281 521 513 301 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=57410 $D=0
M2282 522 514 302 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=62040 $D=0
M2283 523 515 303 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=66670 $D=0
M2284 11 520 1298 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=52780 $D=0
M2285 11 521 1299 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=57410 $D=0
M2286 11 522 1300 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=62040 $D=0
M2287 11 523 1301 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=66670 $D=0
M2288 524 1298 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=52780 $D=0
M2289 525 1299 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=57410 $D=0
M2290 526 1300 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=62040 $D=0
M2291 527 1301 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=66670 $D=0
M2292 520 53 524 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=52780 $D=0
M2293 521 53 525 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=57410 $D=0
M2294 522 53 526 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=62040 $D=0
M2295 523 53 527 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=66670 $D=0
M2296 524 516 320 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=52780 $D=0
M2297 525 517 321 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=57410 $D=0
M2298 526 518 322 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=62040 $D=0
M2299 527 519 323 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=66670 $D=0
M2300 328 528 524 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=52780 $D=0
M2301 329 529 525 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=57410 $D=0
M2302 330 530 526 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=62040 $D=0
M2303 331 531 527 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=66670 $D=0
M2304 528 55 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=52780 $D=0
M2305 529 55 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=57410 $D=0
M2306 530 55 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=62040 $D=0
M2307 531 55 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=66670 $D=0
M2308 11 56 532 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=52780 $D=0
M2309 11 56 533 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=57410 $D=0
M2310 11 56 534 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=62040 $D=0
M2311 11 56 535 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=66670 $D=0
M2312 536 57 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=52780 $D=0
M2313 537 57 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=57410 $D=0
M2314 538 57 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=62040 $D=0
M2315 539 57 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=66670 $D=0
M2316 540 532 300 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=52780 $D=0
M2317 541 533 301 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=57410 $D=0
M2318 542 534 302 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=62040 $D=0
M2319 543 535 303 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=66670 $D=0
M2320 11 540 1302 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=52780 $D=0
M2321 11 541 1303 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=57410 $D=0
M2322 11 542 1304 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=62040 $D=0
M2323 11 543 1305 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=66670 $D=0
M2324 544 1302 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=52780 $D=0
M2325 545 1303 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=57410 $D=0
M2326 546 1304 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=62040 $D=0
M2327 547 1305 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=66670 $D=0
M2328 540 56 544 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=52780 $D=0
M2329 541 56 545 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=57410 $D=0
M2330 542 56 546 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=62040 $D=0
M2331 543 56 547 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=66670 $D=0
M2332 544 536 320 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=52780 $D=0
M2333 545 537 321 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=57410 $D=0
M2334 546 538 322 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=62040 $D=0
M2335 547 539 323 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=66670 $D=0
M2336 328 548 544 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=52780 $D=0
M2337 329 549 545 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=57410 $D=0
M2338 330 550 546 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=62040 $D=0
M2339 331 551 547 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=66670 $D=0
M2340 548 58 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=52780 $D=0
M2341 549 58 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=57410 $D=0
M2342 550 58 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=62040 $D=0
M2343 551 58 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=66670 $D=0
M2344 11 59 552 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=52780 $D=0
M2345 11 59 553 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=57410 $D=0
M2346 11 59 554 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=62040 $D=0
M2347 11 59 555 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=66670 $D=0
M2348 556 60 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=52780 $D=0
M2349 557 60 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=57410 $D=0
M2350 558 60 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=62040 $D=0
M2351 559 60 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=66670 $D=0
M2352 560 552 300 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=52780 $D=0
M2353 561 553 301 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=57410 $D=0
M2354 562 554 302 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=62040 $D=0
M2355 563 555 303 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=66670 $D=0
M2356 11 560 1306 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=52780 $D=0
M2357 11 561 1307 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=57410 $D=0
M2358 11 562 1308 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=62040 $D=0
M2359 11 563 1309 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=66670 $D=0
M2360 564 1306 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=52780 $D=0
M2361 565 1307 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=57410 $D=0
M2362 566 1308 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=62040 $D=0
M2363 567 1309 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=66670 $D=0
M2364 560 59 564 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=52780 $D=0
M2365 561 59 565 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=57410 $D=0
M2366 562 59 566 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=62040 $D=0
M2367 563 59 567 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=66670 $D=0
M2368 564 556 320 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=52780 $D=0
M2369 565 557 321 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=57410 $D=0
M2370 566 558 322 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=62040 $D=0
M2371 567 559 323 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=66670 $D=0
M2372 328 568 564 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=52780 $D=0
M2373 329 569 565 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=57410 $D=0
M2374 330 570 566 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=62040 $D=0
M2375 331 571 567 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=66670 $D=0
M2376 568 61 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=52780 $D=0
M2377 569 61 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=57410 $D=0
M2378 570 61 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=62040 $D=0
M2379 571 61 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=66670 $D=0
M2380 11 62 572 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=52780 $D=0
M2381 11 62 573 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=57410 $D=0
M2382 11 62 574 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=62040 $D=0
M2383 11 62 575 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=66670 $D=0
M2384 576 63 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=52780 $D=0
M2385 577 63 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=57410 $D=0
M2386 578 63 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=62040 $D=0
M2387 579 63 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=66670 $D=0
M2388 580 572 300 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=52780 $D=0
M2389 581 573 301 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=57410 $D=0
M2390 582 574 302 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=62040 $D=0
M2391 583 575 303 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=66670 $D=0
M2392 11 580 1310 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=52780 $D=0
M2393 11 581 1311 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=57410 $D=0
M2394 11 582 1312 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=62040 $D=0
M2395 11 583 1313 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=66670 $D=0
M2396 584 1310 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=52780 $D=0
M2397 585 1311 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=57410 $D=0
M2398 586 1312 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=62040 $D=0
M2399 587 1313 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=66670 $D=0
M2400 580 62 584 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=52780 $D=0
M2401 581 62 585 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=57410 $D=0
M2402 582 62 586 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=62040 $D=0
M2403 583 62 587 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=66670 $D=0
M2404 584 576 320 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=52780 $D=0
M2405 585 577 321 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=57410 $D=0
M2406 586 578 322 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=62040 $D=0
M2407 587 579 323 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=66670 $D=0
M2408 328 588 584 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=52780 $D=0
M2409 329 589 585 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=57410 $D=0
M2410 330 590 586 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=62040 $D=0
M2411 331 591 587 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=66670 $D=0
M2412 588 64 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=52780 $D=0
M2413 589 64 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=57410 $D=0
M2414 590 64 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=62040 $D=0
M2415 591 64 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=66670 $D=0
M2416 11 65 592 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=52780 $D=0
M2417 11 65 593 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=57410 $D=0
M2418 11 65 594 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=62040 $D=0
M2419 11 65 595 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=66670 $D=0
M2420 596 66 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=52780 $D=0
M2421 597 66 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=57410 $D=0
M2422 598 66 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=62040 $D=0
M2423 599 66 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=66670 $D=0
M2424 600 592 300 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=52780 $D=0
M2425 601 593 301 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=57410 $D=0
M2426 602 594 302 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=62040 $D=0
M2427 603 595 303 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=66670 $D=0
M2428 11 600 1314 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=52780 $D=0
M2429 11 601 1315 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=57410 $D=0
M2430 11 602 1316 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=62040 $D=0
M2431 11 603 1317 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=66670 $D=0
M2432 604 1314 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=52780 $D=0
M2433 605 1315 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=57410 $D=0
M2434 606 1316 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=62040 $D=0
M2435 607 1317 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=66670 $D=0
M2436 600 65 604 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=52780 $D=0
M2437 601 65 605 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=57410 $D=0
M2438 602 65 606 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=62040 $D=0
M2439 603 65 607 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=66670 $D=0
M2440 604 596 320 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=52780 $D=0
M2441 605 597 321 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=57410 $D=0
M2442 606 598 322 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=62040 $D=0
M2443 607 599 323 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=66670 $D=0
M2444 328 608 604 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=52780 $D=0
M2445 329 609 605 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=57410 $D=0
M2446 330 610 606 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=62040 $D=0
M2447 331 611 607 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=66670 $D=0
M2448 608 67 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=52780 $D=0
M2449 609 67 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=57410 $D=0
M2450 610 67 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=62040 $D=0
M2451 611 67 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=66670 $D=0
M2452 11 68 612 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=52780 $D=0
M2453 11 68 613 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=57410 $D=0
M2454 11 68 614 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=62040 $D=0
M2455 11 68 615 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=66670 $D=0
M2456 616 69 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=52780 $D=0
M2457 617 69 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=57410 $D=0
M2458 618 69 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=62040 $D=0
M2459 619 69 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=66670 $D=0
M2460 620 612 300 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=52780 $D=0
M2461 621 613 301 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=57410 $D=0
M2462 622 614 302 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=62040 $D=0
M2463 623 615 303 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=66670 $D=0
M2464 11 620 1318 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=52780 $D=0
M2465 11 621 1319 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=57410 $D=0
M2466 11 622 1320 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=62040 $D=0
M2467 11 623 1321 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=66670 $D=0
M2468 624 1318 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=52780 $D=0
M2469 625 1319 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=57410 $D=0
M2470 626 1320 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=62040 $D=0
M2471 627 1321 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=66670 $D=0
M2472 620 68 624 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=52780 $D=0
M2473 621 68 625 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=57410 $D=0
M2474 622 68 626 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=62040 $D=0
M2475 623 68 627 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=66670 $D=0
M2476 624 616 320 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=52780 $D=0
M2477 625 617 321 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=57410 $D=0
M2478 626 618 322 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=62040 $D=0
M2479 627 619 323 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=66670 $D=0
M2480 328 628 624 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=52780 $D=0
M2481 329 629 625 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=57410 $D=0
M2482 330 630 626 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=62040 $D=0
M2483 331 631 627 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=66670 $D=0
M2484 628 70 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=52780 $D=0
M2485 629 70 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=57410 $D=0
M2486 630 70 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=62040 $D=0
M2487 631 70 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=66670 $D=0
M2488 11 71 632 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=52780 $D=0
M2489 11 71 633 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=57410 $D=0
M2490 11 71 634 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=62040 $D=0
M2491 11 71 635 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=66670 $D=0
M2492 636 72 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=52780 $D=0
M2493 637 72 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=57410 $D=0
M2494 638 72 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=62040 $D=0
M2495 639 72 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=66670 $D=0
M2496 640 632 300 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=52780 $D=0
M2497 641 633 301 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=57410 $D=0
M2498 642 634 302 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=62040 $D=0
M2499 643 635 303 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=66670 $D=0
M2500 11 640 1322 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=52780 $D=0
M2501 11 641 1323 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=57410 $D=0
M2502 11 642 1324 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=62040 $D=0
M2503 11 643 1325 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=66670 $D=0
M2504 644 1322 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=52780 $D=0
M2505 645 1323 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=57410 $D=0
M2506 646 1324 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=62040 $D=0
M2507 647 1325 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=66670 $D=0
M2508 640 71 644 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=52780 $D=0
M2509 641 71 645 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=57410 $D=0
M2510 642 71 646 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=62040 $D=0
M2511 643 71 647 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=66670 $D=0
M2512 644 636 320 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=52780 $D=0
M2513 645 637 321 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=57410 $D=0
M2514 646 638 322 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=62040 $D=0
M2515 647 639 323 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=66670 $D=0
M2516 328 648 644 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=52780 $D=0
M2517 329 649 645 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=57410 $D=0
M2518 330 650 646 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=62040 $D=0
M2519 331 651 647 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=66670 $D=0
M2520 648 73 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=52780 $D=0
M2521 649 73 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=57410 $D=0
M2522 650 73 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=62040 $D=0
M2523 651 73 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=66670 $D=0
M2524 11 74 652 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=52780 $D=0
M2525 11 74 653 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=57410 $D=0
M2526 11 74 654 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=62040 $D=0
M2527 11 74 655 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=66670 $D=0
M2528 656 75 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=52780 $D=0
M2529 657 75 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=57410 $D=0
M2530 658 75 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=62040 $D=0
M2531 659 75 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=66670 $D=0
M2532 660 652 300 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=52780 $D=0
M2533 661 653 301 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=57410 $D=0
M2534 662 654 302 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=62040 $D=0
M2535 663 655 303 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=66670 $D=0
M2536 11 660 1326 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=52780 $D=0
M2537 11 661 1327 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=57410 $D=0
M2538 11 662 1328 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=62040 $D=0
M2539 11 663 1329 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=66670 $D=0
M2540 664 1326 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=52780 $D=0
M2541 665 1327 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=57410 $D=0
M2542 666 1328 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=62040 $D=0
M2543 667 1329 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=66670 $D=0
M2544 660 74 664 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=52780 $D=0
M2545 661 74 665 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=57410 $D=0
M2546 662 74 666 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=62040 $D=0
M2547 663 74 667 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=66670 $D=0
M2548 664 656 320 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=52780 $D=0
M2549 665 657 321 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=57410 $D=0
M2550 666 658 322 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=62040 $D=0
M2551 667 659 323 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=66670 $D=0
M2552 328 668 664 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=52780 $D=0
M2553 329 669 665 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=57410 $D=0
M2554 330 670 666 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=62040 $D=0
M2555 331 671 667 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=66670 $D=0
M2556 668 76 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=52780 $D=0
M2557 669 76 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=57410 $D=0
M2558 670 76 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=62040 $D=0
M2559 671 76 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=66670 $D=0
M2560 11 77 672 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=52780 $D=0
M2561 11 77 673 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=57410 $D=0
M2562 11 77 674 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=62040 $D=0
M2563 11 77 675 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=66670 $D=0
M2564 676 78 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=52780 $D=0
M2565 677 78 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=57410 $D=0
M2566 678 78 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=62040 $D=0
M2567 679 78 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=66670 $D=0
M2568 680 672 300 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=52780 $D=0
M2569 681 673 301 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=57410 $D=0
M2570 682 674 302 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=62040 $D=0
M2571 683 675 303 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=66670 $D=0
M2572 11 680 1330 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=52780 $D=0
M2573 11 681 1331 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=57410 $D=0
M2574 11 682 1332 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=62040 $D=0
M2575 11 683 1333 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=66670 $D=0
M2576 684 1330 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=52780 $D=0
M2577 685 1331 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=57410 $D=0
M2578 686 1332 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=62040 $D=0
M2579 687 1333 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=66670 $D=0
M2580 680 77 684 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=52780 $D=0
M2581 681 77 685 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=57410 $D=0
M2582 682 77 686 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=62040 $D=0
M2583 683 77 687 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=66670 $D=0
M2584 684 676 320 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=52780 $D=0
M2585 685 677 321 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=57410 $D=0
M2586 686 678 322 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=62040 $D=0
M2587 687 679 323 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=66670 $D=0
M2588 328 688 684 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=52780 $D=0
M2589 329 689 685 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=57410 $D=0
M2590 330 690 686 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=62040 $D=0
M2591 331 691 687 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=66670 $D=0
M2592 688 79 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=52780 $D=0
M2593 689 79 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=57410 $D=0
M2594 690 79 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=62040 $D=0
M2595 691 79 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=66670 $D=0
M2596 11 80 692 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=52780 $D=0
M2597 11 80 693 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=57410 $D=0
M2598 11 80 694 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=62040 $D=0
M2599 11 80 695 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=66670 $D=0
M2600 696 81 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=52780 $D=0
M2601 697 81 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=57410 $D=0
M2602 698 81 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=62040 $D=0
M2603 699 81 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=66670 $D=0
M2604 700 692 300 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=52780 $D=0
M2605 701 693 301 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=57410 $D=0
M2606 702 694 302 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=62040 $D=0
M2607 703 695 303 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=66670 $D=0
M2608 11 700 1334 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=52780 $D=0
M2609 11 701 1335 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=57410 $D=0
M2610 11 702 1336 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=62040 $D=0
M2611 11 703 1337 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=66670 $D=0
M2612 704 1334 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=52780 $D=0
M2613 705 1335 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=57410 $D=0
M2614 706 1336 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=62040 $D=0
M2615 707 1337 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=66670 $D=0
M2616 700 80 704 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=52780 $D=0
M2617 701 80 705 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=57410 $D=0
M2618 702 80 706 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=62040 $D=0
M2619 703 80 707 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=66670 $D=0
M2620 704 696 320 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=52780 $D=0
M2621 705 697 321 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=57410 $D=0
M2622 706 698 322 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=62040 $D=0
M2623 707 699 323 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=66670 $D=0
M2624 328 708 704 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=52780 $D=0
M2625 329 709 705 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=57410 $D=0
M2626 330 710 706 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=62040 $D=0
M2627 331 711 707 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=66670 $D=0
M2628 708 82 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=52780 $D=0
M2629 709 82 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=57410 $D=0
M2630 710 82 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=62040 $D=0
M2631 711 82 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=66670 $D=0
M2632 11 83 712 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=52780 $D=0
M2633 11 83 713 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=57410 $D=0
M2634 11 83 714 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=62040 $D=0
M2635 11 83 715 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=66670 $D=0
M2636 716 84 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=52780 $D=0
M2637 717 84 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=57410 $D=0
M2638 718 84 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=62040 $D=0
M2639 719 84 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=66670 $D=0
M2640 720 712 300 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=52780 $D=0
M2641 721 713 301 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=57410 $D=0
M2642 722 714 302 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=62040 $D=0
M2643 723 715 303 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=66670 $D=0
M2644 11 720 1338 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=52780 $D=0
M2645 11 721 1339 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=57410 $D=0
M2646 11 722 1340 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=62040 $D=0
M2647 11 723 1341 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=66670 $D=0
M2648 724 1338 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=52780 $D=0
M2649 725 1339 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=57410 $D=0
M2650 726 1340 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=62040 $D=0
M2651 727 1341 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=66670 $D=0
M2652 720 83 724 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=52780 $D=0
M2653 721 83 725 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=57410 $D=0
M2654 722 83 726 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=62040 $D=0
M2655 723 83 727 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=66670 $D=0
M2656 724 716 320 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=52780 $D=0
M2657 725 717 321 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=57410 $D=0
M2658 726 718 322 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=62040 $D=0
M2659 727 719 323 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=66670 $D=0
M2660 328 728 724 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=52780 $D=0
M2661 329 729 725 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=57410 $D=0
M2662 330 730 726 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=62040 $D=0
M2663 331 731 727 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=66670 $D=0
M2664 728 85 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=52780 $D=0
M2665 729 85 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=57410 $D=0
M2666 730 85 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=62040 $D=0
M2667 731 85 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=66670 $D=0
M2668 11 86 732 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=52780 $D=0
M2669 11 86 733 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=57410 $D=0
M2670 11 86 734 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=62040 $D=0
M2671 11 86 735 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=66670 $D=0
M2672 736 87 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=52780 $D=0
M2673 737 87 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=57410 $D=0
M2674 738 87 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=62040 $D=0
M2675 739 87 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=66670 $D=0
M2676 740 732 300 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=52780 $D=0
M2677 741 733 301 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=57410 $D=0
M2678 742 734 302 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=62040 $D=0
M2679 743 735 303 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=66670 $D=0
M2680 11 740 1342 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=52780 $D=0
M2681 11 741 1343 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=57410 $D=0
M2682 11 742 1344 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=62040 $D=0
M2683 11 743 1345 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=66670 $D=0
M2684 744 1342 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=52780 $D=0
M2685 745 1343 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=57410 $D=0
M2686 746 1344 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=62040 $D=0
M2687 747 1345 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=66670 $D=0
M2688 740 86 744 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=52780 $D=0
M2689 741 86 745 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=57410 $D=0
M2690 742 86 746 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=62040 $D=0
M2691 743 86 747 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=66670 $D=0
M2692 744 736 320 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=52780 $D=0
M2693 745 737 321 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=57410 $D=0
M2694 746 738 322 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=62040 $D=0
M2695 747 739 323 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=66670 $D=0
M2696 328 748 744 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=52780 $D=0
M2697 329 749 745 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=57410 $D=0
M2698 330 750 746 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=62040 $D=0
M2699 331 751 747 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=66670 $D=0
M2700 748 88 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=52780 $D=0
M2701 749 88 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=57410 $D=0
M2702 750 88 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=62040 $D=0
M2703 751 88 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=66670 $D=0
M2704 11 89 752 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=52780 $D=0
M2705 11 89 753 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=57410 $D=0
M2706 11 89 754 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=62040 $D=0
M2707 11 89 755 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=66670 $D=0
M2708 756 90 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=52780 $D=0
M2709 757 90 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=57410 $D=0
M2710 758 90 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=62040 $D=0
M2711 759 90 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=66670 $D=0
M2712 760 752 300 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=52780 $D=0
M2713 761 753 301 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=57410 $D=0
M2714 762 754 302 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=62040 $D=0
M2715 763 755 303 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=66670 $D=0
M2716 11 760 1346 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=52780 $D=0
M2717 11 761 1347 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=57410 $D=0
M2718 11 762 1348 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=62040 $D=0
M2719 11 763 1349 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=66670 $D=0
M2720 764 1346 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=52780 $D=0
M2721 765 1347 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=57410 $D=0
M2722 766 1348 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=62040 $D=0
M2723 767 1349 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=66670 $D=0
M2724 760 89 764 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=52780 $D=0
M2725 761 89 765 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=57410 $D=0
M2726 762 89 766 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=62040 $D=0
M2727 763 89 767 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=66670 $D=0
M2728 764 756 320 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=52780 $D=0
M2729 765 757 321 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=57410 $D=0
M2730 766 758 322 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=62040 $D=0
M2731 767 759 323 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=66670 $D=0
M2732 328 768 764 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=52780 $D=0
M2733 329 769 765 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=57410 $D=0
M2734 330 770 766 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=62040 $D=0
M2735 331 771 767 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=66670 $D=0
M2736 768 91 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=52780 $D=0
M2737 769 91 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=57410 $D=0
M2738 770 91 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=62040 $D=0
M2739 771 91 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=66670 $D=0
M2740 11 92 772 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=52780 $D=0
M2741 11 92 773 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=57410 $D=0
M2742 11 92 774 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=62040 $D=0
M2743 11 92 775 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=66670 $D=0
M2744 776 93 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=52780 $D=0
M2745 777 93 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=57410 $D=0
M2746 778 93 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=62040 $D=0
M2747 779 93 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=66670 $D=0
M2748 780 772 300 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=52780 $D=0
M2749 781 773 301 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=57410 $D=0
M2750 782 774 302 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=62040 $D=0
M2751 783 775 303 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=66670 $D=0
M2752 11 780 1350 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=52780 $D=0
M2753 11 781 1351 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=57410 $D=0
M2754 11 782 1352 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=62040 $D=0
M2755 11 783 1353 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=66670 $D=0
M2756 784 1350 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=52780 $D=0
M2757 785 1351 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=57410 $D=0
M2758 786 1352 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=62040 $D=0
M2759 787 1353 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=66670 $D=0
M2760 780 92 784 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=52780 $D=0
M2761 781 92 785 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=57410 $D=0
M2762 782 92 786 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=62040 $D=0
M2763 783 92 787 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=66670 $D=0
M2764 784 776 320 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=52780 $D=0
M2765 785 777 321 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=57410 $D=0
M2766 786 778 322 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=62040 $D=0
M2767 787 779 323 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=66670 $D=0
M2768 328 788 784 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=52780 $D=0
M2769 329 789 785 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=57410 $D=0
M2770 330 790 786 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=62040 $D=0
M2771 331 791 787 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=66670 $D=0
M2772 788 94 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=52780 $D=0
M2773 789 94 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=57410 $D=0
M2774 790 94 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=62040 $D=0
M2775 791 94 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=66670 $D=0
M2776 11 95 792 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=52780 $D=0
M2777 11 95 793 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=57410 $D=0
M2778 11 95 794 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=62040 $D=0
M2779 11 95 795 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=66670 $D=0
M2780 796 96 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=52780 $D=0
M2781 797 96 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=57410 $D=0
M2782 798 96 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=62040 $D=0
M2783 799 96 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=66670 $D=0
M2784 800 792 300 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=52780 $D=0
M2785 801 793 301 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=57410 $D=0
M2786 802 794 302 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=62040 $D=0
M2787 803 795 303 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=66670 $D=0
M2788 11 800 1354 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=52780 $D=0
M2789 11 801 1355 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=57410 $D=0
M2790 11 802 1356 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=62040 $D=0
M2791 11 803 1357 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=66670 $D=0
M2792 804 1354 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=52780 $D=0
M2793 805 1355 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=57410 $D=0
M2794 806 1356 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=62040 $D=0
M2795 807 1357 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=66670 $D=0
M2796 800 95 804 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=52780 $D=0
M2797 801 95 805 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=57410 $D=0
M2798 802 95 806 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=62040 $D=0
M2799 803 95 807 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=66670 $D=0
M2800 804 796 320 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=52780 $D=0
M2801 805 797 321 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=57410 $D=0
M2802 806 798 322 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=62040 $D=0
M2803 807 799 323 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=66670 $D=0
M2804 328 808 804 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=52780 $D=0
M2805 329 809 805 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=57410 $D=0
M2806 330 810 806 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=62040 $D=0
M2807 331 811 807 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=66670 $D=0
M2808 808 97 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=52780 $D=0
M2809 809 97 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=57410 $D=0
M2810 810 97 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=62040 $D=0
M2811 811 97 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=66670 $D=0
M2812 11 98 812 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=52780 $D=0
M2813 11 98 813 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=57410 $D=0
M2814 11 98 814 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=62040 $D=0
M2815 11 98 815 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=66670 $D=0
M2816 816 99 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=52780 $D=0
M2817 817 99 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=57410 $D=0
M2818 818 99 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=62040 $D=0
M2819 819 99 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=66670 $D=0
M2820 820 812 300 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=52780 $D=0
M2821 821 813 301 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=57410 $D=0
M2822 822 814 302 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=62040 $D=0
M2823 823 815 303 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=66670 $D=0
M2824 11 820 1358 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=52780 $D=0
M2825 11 821 1359 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=57410 $D=0
M2826 11 822 1360 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=62040 $D=0
M2827 11 823 1361 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=66670 $D=0
M2828 824 1358 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=52780 $D=0
M2829 825 1359 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=57410 $D=0
M2830 826 1360 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=62040 $D=0
M2831 827 1361 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=66670 $D=0
M2832 820 98 824 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=52780 $D=0
M2833 821 98 825 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=57410 $D=0
M2834 822 98 826 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=62040 $D=0
M2835 823 98 827 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=66670 $D=0
M2836 824 816 320 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=52780 $D=0
M2837 825 817 321 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=57410 $D=0
M2838 826 818 322 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=62040 $D=0
M2839 827 819 323 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=66670 $D=0
M2840 328 828 824 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=52780 $D=0
M2841 329 829 825 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=57410 $D=0
M2842 330 830 826 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=62040 $D=0
M2843 331 831 827 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=66670 $D=0
M2844 828 100 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=52780 $D=0
M2845 829 100 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=57410 $D=0
M2846 830 100 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=62040 $D=0
M2847 831 100 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=66670 $D=0
M2848 11 101 832 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=52780 $D=0
M2849 11 101 833 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=57410 $D=0
M2850 11 101 834 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=62040 $D=0
M2851 11 101 835 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=66670 $D=0
M2852 836 102 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=52780 $D=0
M2853 837 102 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=57410 $D=0
M2854 838 102 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=62040 $D=0
M2855 839 102 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=66670 $D=0
M2856 840 832 300 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=52780 $D=0
M2857 841 833 301 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=57410 $D=0
M2858 842 834 302 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=62040 $D=0
M2859 843 835 303 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=66670 $D=0
M2860 11 840 1362 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=52780 $D=0
M2861 11 841 1363 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=57410 $D=0
M2862 11 842 1364 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=62040 $D=0
M2863 11 843 1365 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=66670 $D=0
M2864 844 1362 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=52780 $D=0
M2865 845 1363 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=57410 $D=0
M2866 846 1364 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=62040 $D=0
M2867 847 1365 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=66670 $D=0
M2868 840 101 844 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=52780 $D=0
M2869 841 101 845 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=57410 $D=0
M2870 842 101 846 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=62040 $D=0
M2871 843 101 847 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=66670 $D=0
M2872 844 836 320 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=52780 $D=0
M2873 845 837 321 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=57410 $D=0
M2874 846 838 322 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=62040 $D=0
M2875 847 839 323 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=66670 $D=0
M2876 328 848 844 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=52780 $D=0
M2877 329 849 845 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=57410 $D=0
M2878 330 850 846 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=62040 $D=0
M2879 331 851 847 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=66670 $D=0
M2880 848 103 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=52780 $D=0
M2881 849 103 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=57410 $D=0
M2882 850 103 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=62040 $D=0
M2883 851 103 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=66670 $D=0
M2884 11 104 852 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=52780 $D=0
M2885 11 104 853 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=57410 $D=0
M2886 11 104 854 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=62040 $D=0
M2887 11 104 855 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=66670 $D=0
M2888 856 105 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=52780 $D=0
M2889 857 105 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=57410 $D=0
M2890 858 105 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=62040 $D=0
M2891 859 105 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=66670 $D=0
M2892 860 852 300 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=52780 $D=0
M2893 861 853 301 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=57410 $D=0
M2894 862 854 302 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=62040 $D=0
M2895 863 855 303 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=66670 $D=0
M2896 11 860 1366 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=52780 $D=0
M2897 11 861 1367 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=57410 $D=0
M2898 11 862 1368 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=62040 $D=0
M2899 11 863 1369 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=66670 $D=0
M2900 864 1366 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=52780 $D=0
M2901 865 1367 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=57410 $D=0
M2902 866 1368 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=62040 $D=0
M2903 867 1369 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=66670 $D=0
M2904 860 104 864 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=52780 $D=0
M2905 861 104 865 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=57410 $D=0
M2906 862 104 866 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=62040 $D=0
M2907 863 104 867 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=66670 $D=0
M2908 864 856 320 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=52780 $D=0
M2909 865 857 321 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=57410 $D=0
M2910 866 858 322 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=62040 $D=0
M2911 867 859 323 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=66670 $D=0
M2912 328 868 864 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=52780 $D=0
M2913 329 869 865 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=57410 $D=0
M2914 330 870 866 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=62040 $D=0
M2915 331 871 867 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=66670 $D=0
M2916 868 106 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=52780 $D=0
M2917 869 106 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=57410 $D=0
M2918 870 106 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=62040 $D=0
M2919 871 106 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=66670 $D=0
M2920 11 107 872 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=52780 $D=0
M2921 11 107 873 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=57410 $D=0
M2922 11 107 874 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=62040 $D=0
M2923 11 107 875 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=66670 $D=0
M2924 876 108 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=52780 $D=0
M2925 877 108 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=57410 $D=0
M2926 878 108 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=62040 $D=0
M2927 879 108 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=66670 $D=0
M2928 880 872 300 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=52780 $D=0
M2929 881 873 301 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=57410 $D=0
M2930 882 874 302 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=62040 $D=0
M2931 883 875 303 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=66670 $D=0
M2932 11 880 1370 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=52780 $D=0
M2933 11 881 1371 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=57410 $D=0
M2934 11 882 1372 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=62040 $D=0
M2935 11 883 1373 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=66670 $D=0
M2936 884 1370 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=52780 $D=0
M2937 885 1371 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=57410 $D=0
M2938 886 1372 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=62040 $D=0
M2939 887 1373 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=66670 $D=0
M2940 880 107 884 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=52780 $D=0
M2941 881 107 885 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=57410 $D=0
M2942 882 107 886 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=62040 $D=0
M2943 883 107 887 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=66670 $D=0
M2944 884 876 320 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=52780 $D=0
M2945 885 877 321 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=57410 $D=0
M2946 886 878 322 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=62040 $D=0
M2947 887 879 323 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=66670 $D=0
M2948 328 888 884 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=52780 $D=0
M2949 329 889 885 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=57410 $D=0
M2950 330 890 886 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=62040 $D=0
M2951 331 891 887 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=66670 $D=0
M2952 888 109 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=52780 $D=0
M2953 889 109 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=57410 $D=0
M2954 890 109 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=62040 $D=0
M2955 891 109 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=66670 $D=0
M2956 11 110 892 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=52780 $D=0
M2957 11 110 893 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=57410 $D=0
M2958 11 110 894 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=62040 $D=0
M2959 11 110 895 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=66670 $D=0
M2960 896 111 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=52780 $D=0
M2961 897 111 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=57410 $D=0
M2962 898 111 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=62040 $D=0
M2963 899 111 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=66670 $D=0
M2964 900 892 300 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=52780 $D=0
M2965 901 893 301 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=57410 $D=0
M2966 902 894 302 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=62040 $D=0
M2967 903 895 303 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=66670 $D=0
M2968 11 900 1374 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=52780 $D=0
M2969 11 901 1375 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=57410 $D=0
M2970 11 902 1376 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=62040 $D=0
M2971 11 903 1377 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=66670 $D=0
M2972 904 1374 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=52780 $D=0
M2973 905 1375 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=57410 $D=0
M2974 906 1376 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=62040 $D=0
M2975 907 1377 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=66670 $D=0
M2976 900 110 904 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=52780 $D=0
M2977 901 110 905 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=57410 $D=0
M2978 902 110 906 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=62040 $D=0
M2979 903 110 907 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=66670 $D=0
M2980 904 896 320 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=52780 $D=0
M2981 905 897 321 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=57410 $D=0
M2982 906 898 322 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=62040 $D=0
M2983 907 899 323 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=66670 $D=0
M2984 328 908 904 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=52780 $D=0
M2985 329 909 905 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=57410 $D=0
M2986 330 910 906 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=62040 $D=0
M2987 331 911 907 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=66670 $D=0
M2988 908 114 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=52780 $D=0
M2989 909 114 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=57410 $D=0
M2990 910 114 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=62040 $D=0
M2991 911 114 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=66670 $D=0
M2992 11 115 912 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=52780 $D=0
M2993 11 115 913 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=57410 $D=0
M2994 11 115 914 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=62040 $D=0
M2995 11 115 915 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=66670 $D=0
M2996 916 116 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=52780 $D=0
M2997 917 116 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=57410 $D=0
M2998 918 116 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=62040 $D=0
M2999 919 116 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=66670 $D=0
M3000 920 912 300 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=52780 $D=0
M3001 921 913 301 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=57410 $D=0
M3002 922 914 302 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=62040 $D=0
M3003 923 915 303 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=66670 $D=0
M3004 11 920 1378 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=52780 $D=0
M3005 11 921 1379 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=57410 $D=0
M3006 11 922 1380 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=62040 $D=0
M3007 11 923 1381 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=66670 $D=0
M3008 924 1378 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=52780 $D=0
M3009 925 1379 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=57410 $D=0
M3010 926 1380 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=62040 $D=0
M3011 927 1381 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=66670 $D=0
M3012 920 115 924 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=52780 $D=0
M3013 921 115 925 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=57410 $D=0
M3014 922 115 926 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=62040 $D=0
M3015 923 115 927 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=66670 $D=0
M3016 924 916 320 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=52780 $D=0
M3017 925 917 321 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=57410 $D=0
M3018 926 918 322 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=62040 $D=0
M3019 927 919 323 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=66670 $D=0
M3020 328 928 924 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=52780 $D=0
M3021 329 929 925 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=57410 $D=0
M3022 330 930 926 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=62040 $D=0
M3023 331 931 927 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=66670 $D=0
M3024 928 120 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=52780 $D=0
M3025 929 120 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=57410 $D=0
M3026 930 120 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=62040 $D=0
M3027 931 120 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=66670 $D=0
M3028 11 121 932 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=52780 $D=0
M3029 11 121 933 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=57410 $D=0
M3030 11 121 934 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=62040 $D=0
M3031 11 121 935 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=66670 $D=0
M3032 936 122 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=52780 $D=0
M3033 937 122 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=57410 $D=0
M3034 938 122 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=62040 $D=0
M3035 939 122 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=66670 $D=0
M3036 8 936 320 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=52780 $D=0
M3037 8 937 321 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=57410 $D=0
M3038 8 938 322 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=62040 $D=0
M3039 8 939 323 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=66670 $D=0
M3040 328 932 8 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=52780 $D=0
M3041 329 933 8 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=57410 $D=0
M3042 330 934 8 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=62040 $D=0
M3043 331 935 8 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=66670 $D=0
M3044 11 944 940 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=52780 $D=0
M3045 11 945 941 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=57410 $D=0
M3046 11 946 942 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=62040 $D=0
M3047 11 947 943 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=66670 $D=0
M3048 944 124 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=52780 $D=0
M3049 945 124 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=57410 $D=0
M3050 946 124 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=62040 $D=0
M3051 947 124 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=66670 $D=0
M3052 1382 320 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=52780 $D=0
M3053 1383 321 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=57410 $D=0
M3054 1384 322 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=62040 $D=0
M3055 1385 323 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=66670 $D=0
M3056 948 944 1382 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=52780 $D=0
M3057 949 945 1383 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=57410 $D=0
M3058 950 946 1384 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=62040 $D=0
M3059 951 947 1385 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=66670 $D=0
M3060 11 948 952 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=52780 $D=0
M3061 11 949 953 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=57410 $D=0
M3062 11 950 954 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=62040 $D=0
M3063 11 951 955 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=66670 $D=0
M3064 1386 952 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=52780 $D=0
M3065 1387 953 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=57410 $D=0
M3066 1388 954 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=62040 $D=0
M3067 1389 955 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=66670 $D=0
M3068 948 940 1386 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=52780 $D=0
M3069 949 941 1387 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=57410 $D=0
M3070 950 942 1388 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=62040 $D=0
M3071 951 943 1389 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=66670 $D=0
M3072 11 960 956 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=52780 $D=0
M3073 11 961 957 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=57410 $D=0
M3074 11 962 958 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=62040 $D=0
M3075 11 963 959 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=66670 $D=0
M3076 960 124 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=52780 $D=0
M3077 961 124 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=57410 $D=0
M3078 962 124 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=62040 $D=0
M3079 963 124 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=66670 $D=0
M3080 1390 328 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=52780 $D=0
M3081 1391 329 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=57410 $D=0
M3082 1392 330 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=62040 $D=0
M3083 1393 331 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=66670 $D=0
M3084 964 960 1390 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=52780 $D=0
M3085 965 961 1391 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=57410 $D=0
M3086 966 962 1392 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=62040 $D=0
M3087 967 963 1393 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=66670 $D=0
M3088 11 964 128 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=52780 $D=0
M3089 11 965 129 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=57410 $D=0
M3090 11 966 130 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=62040 $D=0
M3091 11 967 131 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=66670 $D=0
M3092 1394 128 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=52780 $D=0
M3093 1395 129 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=57410 $D=0
M3094 1396 130 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=62040 $D=0
M3095 1397 131 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=66670 $D=0
M3096 964 956 1394 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=52780 $D=0
M3097 965 957 1395 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=57410 $D=0
M3098 966 958 1396 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=62040 $D=0
M3099 967 959 1397 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=66670 $D=0
M3100 968 132 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=52780 $D=0
M3101 969 132 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=57410 $D=0
M3102 970 132 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=62040 $D=0
M3103 971 132 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=66670 $D=0
M3104 972 132 952 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=52780 $D=0
M3105 973 132 953 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=57410 $D=0
M3106 974 132 954 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=62040 $D=0
M3107 975 132 955 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=66670 $D=0
M3108 133 968 972 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=52780 $D=0
M3109 134 969 973 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=57410 $D=0
M3110 135 970 974 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=62040 $D=0
M3111 136 971 975 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=66670 $D=0
M3112 976 137 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=52780 $D=0
M3113 977 137 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=57410 $D=0
M3114 978 137 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=62040 $D=0
M3115 979 137 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=66670 $D=0
M3116 980 137 128 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=52780 $D=0
M3117 981 137 129 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=57410 $D=0
M3118 982 137 130 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=62040 $D=0
M3119 983 137 131 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=66670 $D=0
M3120 1398 976 980 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=52780 $D=0
M3121 1399 977 981 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=57410 $D=0
M3122 1400 978 982 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=62040 $D=0
M3123 1401 979 983 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=66670 $D=0
M3124 11 128 1398 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=52780 $D=0
M3125 11 129 1399 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=57410 $D=0
M3126 11 130 1400 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=62040 $D=0
M3127 11 131 1401 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=66670 $D=0
M3128 984 138 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=52780 $D=0
M3129 985 138 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=57410 $D=0
M3130 986 138 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=62040 $D=0
M3131 987 138 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=66670 $D=0
M3132 988 138 980 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=52780 $D=0
M3133 989 138 981 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=57410 $D=0
M3134 990 138 982 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=62040 $D=0
M3135 991 138 983 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=66670 $D=0
M3136 13 984 988 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=52780 $D=0
M3137 14 985 989 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=57410 $D=0
M3138 15 986 990 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=62040 $D=0
M3139 16 987 991 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=66670 $D=0
M3140 995 992 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=52780 $D=0
M3141 996 993 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=57410 $D=0
M3142 997 994 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=62040 $D=0
M3143 998 139 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=66670 $D=0
M3144 11 1003 999 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=52780 $D=0
M3145 11 1004 1000 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=57410 $D=0
M3146 11 1005 1001 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=62040 $D=0
M3147 11 1006 1002 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=66670 $D=0
M3148 1007 972 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=52780 $D=0
M3149 1008 973 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=57410 $D=0
M3150 1009 974 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=62040 $D=0
M3151 1010 975 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=66670 $D=0
M3152 1003 972 992 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=52780 $D=0
M3153 1004 973 993 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=57410 $D=0
M3154 1005 974 994 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=62040 $D=0
M3155 1006 975 139 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=66670 $D=0
M3156 995 1007 1003 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=52780 $D=0
M3157 996 1008 1004 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=57410 $D=0
M3158 997 1009 1005 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=62040 $D=0
M3159 998 1010 1006 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=66670 $D=0
M3160 1011 999 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=52780 $D=0
M3161 1012 1000 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=57410 $D=0
M3162 1013 1001 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=62040 $D=0
M3163 1014 1002 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=66670 $D=0
M3164 140 999 988 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=52780 $D=0
M3165 992 1000 989 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=57410 $D=0
M3166 993 1001 990 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=62040 $D=0
M3167 994 1002 991 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=66670 $D=0
M3168 972 1011 140 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=52780 $D=0
M3169 973 1012 992 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=57410 $D=0
M3170 974 1013 993 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=62040 $D=0
M3171 975 1014 994 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=66670 $D=0
M3172 1015 140 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=52780 $D=0
M3173 1016 992 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=57410 $D=0
M3174 1017 993 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=62040 $D=0
M3175 1018 994 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=66670 $D=0
M3176 1019 999 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=52780 $D=0
M3177 1020 1000 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=57410 $D=0
M3178 1021 1001 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=62040 $D=0
M3179 1022 1002 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=66670 $D=0
M3180 1023 999 1015 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=52780 $D=0
M3181 1024 1000 1016 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=57410 $D=0
M3182 1025 1001 1017 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=62040 $D=0
M3183 1026 1002 1018 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=66670 $D=0
M3184 988 1019 1023 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=52780 $D=0
M3185 989 1020 1024 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=57410 $D=0
M3186 990 1021 1025 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=62040 $D=0
M3187 991 1022 1026 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=66670 $D=0
M3188 1422 972 11 11 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=52420 $D=0
M3189 1423 973 11 11 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=57050 $D=0
M3190 1424 974 11 11 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=61680 $D=0
M3191 1425 975 11 11 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=66310 $D=0
M3192 1027 988 1422 11 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=52420 $D=0
M3193 1028 989 1423 11 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=57050 $D=0
M3194 1029 990 1424 11 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=61680 $D=0
M3195 1030 991 1425 11 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=66310 $D=0
M3196 1031 1023 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=52780 $D=0
M3197 1032 1024 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=57410 $D=0
M3198 1033 1025 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=62040 $D=0
M3199 1034 1026 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=66670 $D=0
M3200 1035 972 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=52780 $D=0
M3201 1036 973 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=57410 $D=0
M3202 1037 974 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=62040 $D=0
M3203 1038 975 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=66670 $D=0
M3204 11 988 1035 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=52780 $D=0
M3205 11 989 1036 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=57410 $D=0
M3206 11 990 1037 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=62040 $D=0
M3207 11 991 1038 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=66670 $D=0
M3208 1039 972 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=52780 $D=0
M3209 1040 973 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=57410 $D=0
M3210 1041 974 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=62040 $D=0
M3211 1042 975 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=66670 $D=0
M3212 11 988 1039 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=52780 $D=0
M3213 11 989 1040 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=57410 $D=0
M3214 11 990 1041 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=62040 $D=0
M3215 11 991 1042 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=66670 $D=0
M3216 1426 972 11 11 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=52600 $D=0
M3217 1427 973 11 11 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=57230 $D=0
M3218 1428 974 11 11 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=61860 $D=0
M3219 1429 975 11 11 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=66490 $D=0
M3220 1047 988 1426 11 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=52600 $D=0
M3221 1048 989 1427 11 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=57230 $D=0
M3222 1049 990 1428 11 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=61860 $D=0
M3223 1050 991 1429 11 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=66490 $D=0
M3224 11 1039 1047 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=52780 $D=0
M3225 11 1040 1048 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=57410 $D=0
M3226 11 1041 1049 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=62040 $D=0
M3227 11 1042 1050 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=66670 $D=0
M3228 1051 144 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=52780 $D=0
M3229 1052 144 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=57410 $D=0
M3230 1053 144 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=62040 $D=0
M3231 1054 144 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=66670 $D=0
M3232 1055 144 1027 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=52780 $D=0
M3233 1056 144 1028 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=57410 $D=0
M3234 1057 144 1029 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=62040 $D=0
M3235 1058 144 1030 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=66670 $D=0
M3236 1035 1051 1055 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=52780 $D=0
M3237 1036 1052 1056 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=57410 $D=0
M3238 1037 1053 1057 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=62040 $D=0
M3239 1038 1054 1058 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=66670 $D=0
M3240 1059 144 1031 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=52780 $D=0
M3241 1060 144 1032 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=57410 $D=0
M3242 1061 144 1033 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=62040 $D=0
M3243 1062 144 1034 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=66670 $D=0
M3244 1047 1051 1059 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=52780 $D=0
M3245 1048 1052 1060 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=57410 $D=0
M3246 1049 1053 1061 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=62040 $D=0
M3247 1050 1054 1062 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=66670 $D=0
M3248 1063 145 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=52780 $D=0
M3249 1064 145 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=57410 $D=0
M3250 1065 145 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=62040 $D=0
M3251 1066 145 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=66670 $D=0
M3252 1067 145 1059 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=52780 $D=0
M3253 1068 145 1060 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=57410 $D=0
M3254 1069 145 1061 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=62040 $D=0
M3255 1070 145 1062 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=66670 $D=0
M3256 1055 1063 1067 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=52780 $D=0
M3257 1056 1064 1068 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=57410 $D=0
M3258 1057 1065 1069 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=62040 $D=0
M3259 1058 1066 1070 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=66670 $D=0
M3260 17 1067 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=52780 $D=0
M3261 18 1068 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=57410 $D=0
M3262 19 1069 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=62040 $D=0
M3263 20 1070 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=66670 $D=0
M3264 1071 146 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=52780 $D=0
M3265 1072 146 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=57410 $D=0
M3266 1073 146 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=62040 $D=0
M3267 1074 146 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=66670 $D=0
M3268 1077 146 1075 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=52780 $D=0
M3269 1078 146 1076 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=57410 $D=0
M3270 1079 146 147 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=62040 $D=0
M3271 1080 146 148 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=66670 $D=0
M3272 149 1071 1077 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=52780 $D=0
M3273 150 1072 1078 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=57410 $D=0
M3274 1075 1073 1079 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=62040 $D=0
M3275 1076 1074 1080 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=66670 $D=0
M3276 1081 146 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=52780 $D=0
M3277 1082 146 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=57410 $D=0
M3278 1083 146 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=62040 $D=0
M3279 1084 146 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=66670 $D=0
M3280 1085 146 151 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=52780 $D=0
M3281 1086 146 152 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=57410 $D=0
M3282 1087 146 153 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=62040 $D=0
M3283 1088 146 154 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=66670 $D=0
M3284 155 1081 1085 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=52780 $D=0
M3285 156 1082 1086 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=57410 $D=0
M3286 157 1083 1087 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=62040 $D=0
M3287 158 1084 1088 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=66670 $D=0
M3288 1089 146 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=52780 $D=0
M3289 1090 146 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=57410 $D=0
M3290 1091 146 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=62040 $D=0
M3291 1092 146 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=66670 $D=0
M3292 1093 146 141 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=52780 $D=0
M3293 1094 146 143 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=57410 $D=0
M3294 1095 146 142 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=62040 $D=0
M3295 1096 146 159 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=66670 $D=0
M3296 160 1089 1093 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=52780 $D=0
M3297 118 1090 1094 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=57410 $D=0
M3298 119 1091 1095 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=62040 $D=0
M3299 123 1092 1096 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=66670 $D=0
M3300 1097 146 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=52780 $D=0
M3301 1098 146 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=57410 $D=0
M3302 1099 146 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=62040 $D=0
M3303 1100 146 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=66670 $D=0
M3304 1101 146 161 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=52780 $D=0
M3305 1102 146 162 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=57410 $D=0
M3306 1103 146 163 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=62040 $D=0
M3307 1104 146 164 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=66670 $D=0
M3308 165 1097 1101 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=52780 $D=0
M3309 166 1098 1102 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=57410 $D=0
M3310 167 1099 1103 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=62040 $D=0
M3311 168 1100 1104 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=66670 $D=0
M3312 1105 146 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=52780 $D=0
M3313 1106 146 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=57410 $D=0
M3314 1107 146 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=62040 $D=0
M3315 1108 146 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=66670 $D=0
M3316 1109 146 169 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=52780 $D=0
M3317 1110 146 170 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=57410 $D=0
M3318 1111 146 171 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=62040 $D=0
M3319 1112 146 172 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=66670 $D=0
M3320 173 1105 1109 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=52780 $D=0
M3321 173 1106 1110 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=57410 $D=0
M3322 173 1107 1111 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=62040 $D=0
M3323 173 1108 1112 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=66670 $D=0
M3324 11 972 1402 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=52780 $D=0
M3325 11 973 1403 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=57410 $D=0
M3326 11 974 1404 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=62040 $D=0
M3327 11 975 1405 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=66670 $D=0
M3328 150 1402 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=52780 $D=0
M3329 1075 1403 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=57410 $D=0
M3330 1076 1404 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=62040 $D=0
M3331 147 1405 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=66670 $D=0
M3332 1113 174 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=52780 $D=0
M3333 1114 174 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=57410 $D=0
M3334 1115 174 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=62040 $D=0
M3335 1116 174 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=66670 $D=0
M3336 157 174 150 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=52780 $D=0
M3337 158 174 1075 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=57410 $D=0
M3338 151 174 1076 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=62040 $D=0
M3339 152 174 147 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=66670 $D=0
M3340 1077 1113 157 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=52780 $D=0
M3341 1078 1114 158 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=57410 $D=0
M3342 1079 1115 151 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=62040 $D=0
M3343 1080 1116 152 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=66670 $D=0
M3344 1117 175 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=52780 $D=0
M3345 1118 175 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=57410 $D=0
M3346 1119 175 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=62040 $D=0
M3347 1120 175 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=66670 $D=0
M3348 176 175 157 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=52780 $D=0
M3349 125 175 158 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=57410 $D=0
M3350 126 175 151 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=62040 $D=0
M3351 127 175 152 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=66670 $D=0
M3352 1085 1117 176 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=52780 $D=0
M3353 1086 1118 125 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=57410 $D=0
M3354 1087 1119 126 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=62040 $D=0
M3355 1088 1120 127 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=66670 $D=0
M3356 1121 177 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=52780 $D=0
M3357 1122 177 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=57410 $D=0
M3358 1123 177 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=62040 $D=0
M3359 1124 177 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=66670 $D=0
M3360 178 177 176 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=52780 $D=0
M3361 112 177 125 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=57410 $D=0
M3362 113 177 126 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=62040 $D=0
M3363 117 177 127 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=66670 $D=0
M3364 1093 1121 178 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=52780 $D=0
M3365 1094 1122 112 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=57410 $D=0
M3366 1095 1123 113 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=62040 $D=0
M3367 1096 1124 117 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=66670 $D=0
M3368 1125 179 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=52780 $D=0
M3369 1126 179 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=57410 $D=0
M3370 1127 179 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=62040 $D=0
M3371 1128 179 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=66670 $D=0
M3372 180 179 178 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=52780 $D=0
M3373 181 179 112 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=57410 $D=0
M3374 182 179 113 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=62040 $D=0
M3375 183 179 117 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=66670 $D=0
M3376 1101 1125 180 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=52780 $D=0
M3377 1102 1126 181 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=57410 $D=0
M3378 1103 1127 182 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=62040 $D=0
M3379 1104 1128 183 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=66670 $D=0
M3380 1129 184 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=52780 $D=0
M3381 1130 184 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=57410 $D=0
M3382 1131 184 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=62040 $D=0
M3383 1132 184 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=66670 $D=0
M3384 272 184 180 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=52780 $D=0
M3385 273 184 181 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=57410 $D=0
M3386 274 184 182 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=62040 $D=0
M3387 275 184 183 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=66670 $D=0
M3388 1109 1129 272 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=52780 $D=0
M3389 1110 1130 273 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=57410 $D=0
M3390 1111 1131 274 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=62040 $D=0
M3391 1112 1132 275 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=66670 $D=0
M3392 1133 185 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=52780 $D=0
M3393 1134 185 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=57410 $D=0
M3394 1135 185 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=62040 $D=0
M3395 1136 185 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=66670 $D=0
M3396 1137 185 128 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=52780 $D=0
M3397 1138 185 129 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=57410 $D=0
M3398 1139 185 130 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=62040 $D=0
M3399 1140 185 131 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=66670 $D=0
M3400 13 1133 1137 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=52780 $D=0
M3401 14 1134 1138 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=57410 $D=0
M3402 15 1135 1139 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=62040 $D=0
M3403 16 1136 1140 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=66670 $D=0
M3404 1141 952 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=52780 $D=0
M3405 1142 953 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=57410 $D=0
M3406 1143 954 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=62040 $D=0
M3407 1144 955 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=66670 $D=0
M3408 11 1137 1141 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=52780 $D=0
M3409 11 1138 1142 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=57410 $D=0
M3410 11 1139 1143 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=62040 $D=0
M3411 11 1140 1144 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=66670 $D=0
M3412 1430 952 11 11 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=52600 $D=0
M3413 1431 953 11 11 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=57230 $D=0
M3414 1432 954 11 11 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=61860 $D=0
M3415 1433 955 11 11 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=66490 $D=0
M3416 1149 1137 1430 11 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=52600 $D=0
M3417 1150 1138 1431 11 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=57230 $D=0
M3418 1151 1139 1432 11 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=61860 $D=0
M3419 1152 1140 1433 11 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=66490 $D=0
M3420 11 1141 1149 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=52780 $D=0
M3421 11 1142 1150 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=57410 $D=0
M3422 11 1143 1151 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=62040 $D=0
M3423 11 1144 1152 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=66670 $D=0
M3424 1406 186 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=52780 $D=0
M3425 1407 1153 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=57410 $D=0
M3426 1408 1154 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=62040 $D=0
M3427 1409 1155 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=66670 $D=0
M3428 11 1149 1406 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=52780 $D=0
M3429 11 1150 1407 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=57410 $D=0
M3430 11 1151 1408 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=62040 $D=0
M3431 11 1152 1409 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=66670 $D=0
M3432 1153 1406 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=52780 $D=0
M3433 1154 1407 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=57410 $D=0
M3434 1155 1408 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=62040 $D=0
M3435 187 1409 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=66670 $D=0
M3436 1434 952 11 11 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=52420 $D=0
M3437 1435 953 11 11 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=57050 $D=0
M3438 1436 954 11 11 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=61680 $D=0
M3439 1437 955 11 11 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=66310 $D=0
M3440 1156 1160 1434 11 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=52420 $D=0
M3441 1157 1161 1435 11 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=57050 $D=0
M3442 1158 1162 1436 11 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=61680 $D=0
M3443 1159 1163 1437 11 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=66310 $D=0
M3444 1160 1137 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=52780 $D=0
M3445 1161 1138 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=57410 $D=0
M3446 1162 1139 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=62040 $D=0
M3447 1163 1140 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=66670 $D=0
M3448 1164 1156 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=52780 $D=0
M3449 1165 1157 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=57410 $D=0
M3450 1166 1158 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=62040 $D=0
M3451 1167 1159 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=66670 $D=0
M3452 11 186 1164 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=52780 $D=0
M3453 11 1153 1165 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=57410 $D=0
M3454 11 1154 1166 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=62040 $D=0
M3455 11 1155 1167 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=66670 $D=0
M3456 1171 188 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=52780 $D=0
M3457 1172 1168 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=57410 $D=0
M3458 1173 1169 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=62040 $D=0
M3459 1174 1170 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=66670 $D=0
M3460 1168 1164 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=52780 $D=0
M3461 1169 1165 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=57410 $D=0
M3462 1170 1166 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=62040 $D=0
M3463 189 1167 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=66670 $D=0
M3464 11 1171 1168 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=52780 $D=0
M3465 11 1172 1169 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=57410 $D=0
M3466 11 1173 1170 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=62040 $D=0
M3467 11 1174 189 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=66670 $D=0
M3468 1178 1175 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=52780 $D=0
M3469 1179 1176 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=57410 $D=0
M3470 1180 1177 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=62040 $D=0
M3471 1181 190 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=66670 $D=0
M3472 11 1186 1182 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=52780 $D=0
M3473 11 1187 1183 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=57410 $D=0
M3474 11 1188 1184 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=62040 $D=0
M3475 11 1189 1185 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=66670 $D=0
M3476 1190 133 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=52780 $D=0
M3477 1191 134 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=57410 $D=0
M3478 1192 135 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=62040 $D=0
M3479 1193 136 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=66670 $D=0
M3480 1186 133 1175 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=52780 $D=0
M3481 1187 134 1176 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=57410 $D=0
M3482 1188 135 1177 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=62040 $D=0
M3483 1189 136 190 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=66670 $D=0
M3484 1178 1190 1186 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=52780 $D=0
M3485 1179 1191 1187 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=57410 $D=0
M3486 1180 1192 1188 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=62040 $D=0
M3487 1181 1193 1189 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=66670 $D=0
M3488 1194 1182 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=52780 $D=0
M3489 1195 1183 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=57410 $D=0
M3490 1196 1184 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=62040 $D=0
M3491 1197 1185 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=66670 $D=0
M3492 191 1182 8 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=52780 $D=0
M3493 1175 1183 8 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=57410 $D=0
M3494 1176 1184 8 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=62040 $D=0
M3495 1177 1185 8 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=66670 $D=0
M3496 133 1194 191 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=52780 $D=0
M3497 134 1195 1175 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=57410 $D=0
M3498 135 1196 1176 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=62040 $D=0
M3499 136 1197 1177 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=66670 $D=0
M3500 1198 191 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=52780 $D=0
M3501 1199 1175 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=57410 $D=0
M3502 1200 1176 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=62040 $D=0
M3503 1201 1177 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=66670 $D=0
M3504 1202 1182 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=52780 $D=0
M3505 1203 1183 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=57410 $D=0
M3506 1204 1184 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=62040 $D=0
M3507 1205 1185 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=66670 $D=0
M3508 276 1182 1198 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=52780 $D=0
M3509 277 1183 1199 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=57410 $D=0
M3510 278 1184 1200 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=62040 $D=0
M3511 279 1185 1201 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=66670 $D=0
M3512 8 1202 276 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=52780 $D=0
M3513 8 1203 277 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=57410 $D=0
M3514 8 1204 278 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=62040 $D=0
M3515 8 1205 279 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=66670 $D=0
M3516 1206 192 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=52780 $D=0
M3517 1207 192 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=57410 $D=0
M3518 1208 192 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=62040 $D=0
M3519 1209 192 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=66670 $D=0
M3520 1210 192 276 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=52780 $D=0
M3521 1211 192 277 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=57410 $D=0
M3522 1212 192 278 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=62040 $D=0
M3523 1213 192 279 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=66670 $D=0
M3524 17 1206 1210 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=52780 $D=0
M3525 18 1207 1211 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=57410 $D=0
M3526 19 1208 1212 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=62040 $D=0
M3527 20 1209 1213 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=66670 $D=0
M3528 1214 193 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=52780 $D=0
M3529 1215 193 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=57410 $D=0
M3530 1216 193 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=62040 $D=0
M3531 1217 193 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=66670 $D=0
M3532 1218 193 1210 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=52780 $D=0
M3533 1219 193 1211 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=57410 $D=0
M3534 1220 193 1212 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=62040 $D=0
M3535 1221 193 1213 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=66670 $D=0
M3536 8 1214 1218 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=52780 $D=0
M3537 8 1215 1219 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=57410 $D=0
M3538 8 1216 1220 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=62040 $D=0
M3539 8 1217 1221 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=66670 $D=0
M3540 1222 124 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=52780 $D=0
M3541 1223 124 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=57410 $D=0
M3542 1224 124 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=62040 $D=0
M3543 1225 124 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=66670 $D=0
M3544 11 1222 1226 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=52780 $D=0
M3545 11 1223 1227 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=57410 $D=0
M3546 11 1224 1228 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=62040 $D=0
M3547 11 1225 1229 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=66670 $D=0
M3548 1230 124 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=52780 $D=0
M3549 1231 124 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=57410 $D=0
M3550 1232 124 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=62040 $D=0
M3551 1233 124 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=66670 $D=0
M3552 1234 1226 1218 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=52780 $D=0
M3553 1235 1227 1219 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=57410 $D=0
M3554 1236 1228 1220 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=62040 $D=0
M3555 1237 1229 1221 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=66670 $D=0
M3556 11 1234 1410 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=52780 $D=0
M3557 11 1235 1411 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=57410 $D=0
M3558 11 1236 1412 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=62040 $D=0
M3559 11 1237 1413 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=66670 $D=0
M3560 1238 1410 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=52780 $D=0
M3561 1239 1411 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=57410 $D=0
M3562 1240 1412 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=62040 $D=0
M3563 1241 1413 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=66670 $D=0
M3564 1234 1222 1238 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=52780 $D=0
M3565 1235 1223 1239 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=57410 $D=0
M3566 1236 1224 1240 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=62040 $D=0
M3567 1237 1225 1241 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=66670 $D=0
M3568 1242 1230 1238 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=52780 $D=0
M3569 1243 1231 1239 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=57410 $D=0
M3570 1244 1232 1240 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=62040 $D=0
M3571 1245 1233 1241 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=66670 $D=0
M3572 11 1250 1246 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=52780 $D=0
M3573 11 1251 1247 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=57410 $D=0
M3574 11 1252 1248 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=62040 $D=0
M3575 11 1253 1249 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=66670 $D=0
M3576 1250 124 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=52780 $D=0
M3577 1251 124 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=57410 $D=0
M3578 1252 124 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=62040 $D=0
M3579 1253 124 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=66670 $D=0
M3580 1414 1242 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=52780 $D=0
M3581 1415 1243 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=57410 $D=0
M3582 1416 1244 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=62040 $D=0
M3583 1417 1245 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=66670 $D=0
M3584 1254 1250 1414 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=52780 $D=0
M3585 1255 1251 1415 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=57410 $D=0
M3586 1256 1252 1416 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=62040 $D=0
M3587 1257 1253 1417 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=66670 $D=0
M3588 11 1254 133 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=52780 $D=0
M3589 11 1255 134 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=57410 $D=0
M3590 11 1256 135 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=62040 $D=0
M3591 11 1257 136 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=66670 $D=0
M3592 1418 133 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=52780 $D=0
M3593 1419 134 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=57410 $D=0
M3594 1420 135 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=62040 $D=0
M3595 1421 136 11 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=66670 $D=0
M3596 1254 1246 1418 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=52780 $D=0
M3597 1255 1247 1419 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=57410 $D=0
M3598 1256 1248 1420 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=62040 $D=0
M3599 1257 1249 1421 11 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=66670 $D=0
.ENDS
***************************************
.SUBCKT ICV_37 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 108 109 110 111 113 114 115 116 117 119 120 121 122 123
+ 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141 142 143
+ 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162 163
+ 164 165 166 167 168
** N=816 EP=165 IP=1514 FDC=1800
M0 201 1 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=42270 $D=1
M1 202 1 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=46900 $D=1
M2 203 201 2 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=42270 $D=1
M3 204 202 3 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=46900 $D=1
M4 6 1 203 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=42270 $D=1
M5 6 1 204 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=46900 $D=1
M6 205 201 4 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=42270 $D=1
M7 206 202 4 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=46900 $D=1
M8 5 1 205 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=42270 $D=1
M9 5 1 206 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=46900 $D=1
M10 207 201 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=42270 $D=1
M11 208 202 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=46900 $D=1
M12 6 1 207 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=42270 $D=1
M13 6 1 208 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=46900 $D=1
M14 211 209 207 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=42270 $D=1
M15 212 210 208 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=46900 $D=1
M16 209 7 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=42270 $D=1
M17 210 7 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=46900 $D=1
M18 213 209 205 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=42270 $D=1
M19 214 210 206 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=46900 $D=1
M20 203 7 213 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=42270 $D=1
M21 204 7 214 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=46900 $D=1
M22 215 8 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=42270 $D=1
M23 216 8 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=46900 $D=1
M24 217 215 213 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=42270 $D=1
M25 218 216 214 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=46900 $D=1
M26 211 8 217 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=42270 $D=1
M27 212 8 218 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=46900 $D=1
M28 219 10 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=42270 $D=1
M29 220 10 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=46900 $D=1
M30 221 219 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=42270 $D=1
M31 222 220 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=46900 $D=1
M32 11 10 221 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=42270 $D=1
M33 12 10 222 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=46900 $D=1
M34 223 219 13 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=42270 $D=1
M35 224 220 14 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=46900 $D=1
M36 225 10 223 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=42270 $D=1
M37 226 10 224 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=46900 $D=1
M38 229 219 227 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=42270 $D=1
M39 230 220 228 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=46900 $D=1
M40 217 10 229 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=42270 $D=1
M41 218 10 230 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=46900 $D=1
M42 233 231 229 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=42270 $D=1
M43 234 232 230 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=46900 $D=1
M44 231 15 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=42270 $D=1
M45 232 15 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=46900 $D=1
M46 235 231 223 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=42270 $D=1
M47 236 232 224 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=46900 $D=1
M48 221 15 235 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=42270 $D=1
M49 222 15 236 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=46900 $D=1
M50 237 16 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=42270 $D=1
M51 238 16 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=46900 $D=1
M52 239 237 235 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=42270 $D=1
M53 240 238 236 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=46900 $D=1
M54 233 16 239 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=42270 $D=1
M55 234 16 240 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=46900 $D=1
M56 6 17 241 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=42270 $D=1
M57 6 17 242 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=46900 $D=1
M58 243 18 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=42270 $D=1
M59 244 18 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=46900 $D=1
M60 245 17 239 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=42270 $D=1
M61 246 17 240 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=46900 $D=1
M62 6 245 715 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=42270 $D=1
M63 6 246 716 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=46900 $D=1
M64 247 715 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=42270 $D=1
M65 248 716 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=46900 $D=1
M66 245 241 247 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=42270 $D=1
M67 246 242 248 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=46900 $D=1
M68 247 18 249 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=42270 $D=1
M69 248 18 250 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=46900 $D=1
M70 253 19 247 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=42270 $D=1
M71 254 19 248 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=46900 $D=1
M72 251 19 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=42270 $D=1
M73 252 19 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=46900 $D=1
M74 6 20 255 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=42270 $D=1
M75 6 20 256 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=46900 $D=1
M76 257 21 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=42270 $D=1
M77 258 21 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=46900 $D=1
M78 259 20 239 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=42270 $D=1
M79 260 20 240 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=46900 $D=1
M80 6 259 717 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=42270 $D=1
M81 6 260 718 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=46900 $D=1
M82 261 717 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=42270 $D=1
M83 262 718 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=46900 $D=1
M84 259 255 261 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=42270 $D=1
M85 260 256 262 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=46900 $D=1
M86 261 21 249 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=42270 $D=1
M87 262 21 250 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=46900 $D=1
M88 253 22 261 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=42270 $D=1
M89 254 22 262 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=46900 $D=1
M90 263 22 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=42270 $D=1
M91 264 22 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=46900 $D=1
M92 6 23 265 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=42270 $D=1
M93 6 23 266 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=46900 $D=1
M94 267 24 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=42270 $D=1
M95 268 24 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=46900 $D=1
M96 269 23 239 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=42270 $D=1
M97 270 23 240 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=46900 $D=1
M98 6 269 719 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=42270 $D=1
M99 6 270 720 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=46900 $D=1
M100 271 719 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=42270 $D=1
M101 272 720 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=46900 $D=1
M102 269 265 271 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=42270 $D=1
M103 270 266 272 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=46900 $D=1
M104 271 24 249 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=42270 $D=1
M105 272 24 250 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=46900 $D=1
M106 253 25 271 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=42270 $D=1
M107 254 25 272 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=46900 $D=1
M108 273 25 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=42270 $D=1
M109 274 25 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=46900 $D=1
M110 6 26 275 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=42270 $D=1
M111 6 26 276 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=46900 $D=1
M112 277 27 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=42270 $D=1
M113 278 27 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=46900 $D=1
M114 279 26 239 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=42270 $D=1
M115 280 26 240 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=46900 $D=1
M116 6 279 721 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=42270 $D=1
M117 6 280 722 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=46900 $D=1
M118 281 721 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=42270 $D=1
M119 282 722 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=46900 $D=1
M120 279 275 281 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=42270 $D=1
M121 280 276 282 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=46900 $D=1
M122 281 27 249 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=42270 $D=1
M123 282 27 250 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=46900 $D=1
M124 253 28 281 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=42270 $D=1
M125 254 28 282 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=46900 $D=1
M126 283 28 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=42270 $D=1
M127 284 28 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=46900 $D=1
M128 6 29 285 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=42270 $D=1
M129 6 29 286 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=46900 $D=1
M130 287 30 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=42270 $D=1
M131 288 30 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=46900 $D=1
M132 289 29 239 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=42270 $D=1
M133 290 29 240 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=46900 $D=1
M134 6 289 723 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=42270 $D=1
M135 6 290 724 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=46900 $D=1
M136 291 723 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=42270 $D=1
M137 292 724 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=46900 $D=1
M138 289 285 291 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=42270 $D=1
M139 290 286 292 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=46900 $D=1
M140 291 30 249 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=42270 $D=1
M141 292 30 250 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=46900 $D=1
M142 253 31 291 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=42270 $D=1
M143 254 31 292 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=46900 $D=1
M144 293 31 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=42270 $D=1
M145 294 31 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=46900 $D=1
M146 6 32 295 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=42270 $D=1
M147 6 32 296 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=46900 $D=1
M148 297 33 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=42270 $D=1
M149 298 33 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=46900 $D=1
M150 299 32 239 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=42270 $D=1
M151 300 32 240 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=46900 $D=1
M152 6 299 725 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=42270 $D=1
M153 6 300 726 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=46900 $D=1
M154 301 725 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=42270 $D=1
M155 302 726 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=46900 $D=1
M156 299 295 301 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=42270 $D=1
M157 300 296 302 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=46900 $D=1
M158 301 33 249 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=42270 $D=1
M159 302 33 250 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=46900 $D=1
M160 253 34 301 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=42270 $D=1
M161 254 34 302 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=46900 $D=1
M162 303 34 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=42270 $D=1
M163 304 34 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=46900 $D=1
M164 6 35 305 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=42270 $D=1
M165 6 35 306 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=46900 $D=1
M166 307 36 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=42270 $D=1
M167 308 36 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=46900 $D=1
M168 309 35 239 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=42270 $D=1
M169 310 35 240 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=46900 $D=1
M170 6 309 727 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=42270 $D=1
M171 6 310 728 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=46900 $D=1
M172 311 727 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=42270 $D=1
M173 312 728 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=46900 $D=1
M174 309 305 311 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=42270 $D=1
M175 310 306 312 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=46900 $D=1
M176 311 36 249 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=42270 $D=1
M177 312 36 250 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=46900 $D=1
M178 253 37 311 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=42270 $D=1
M179 254 37 312 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=46900 $D=1
M180 313 37 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=42270 $D=1
M181 314 37 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=46900 $D=1
M182 6 38 315 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=42270 $D=1
M183 6 38 316 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=46900 $D=1
M184 317 39 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=42270 $D=1
M185 318 39 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=46900 $D=1
M186 319 38 239 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=42270 $D=1
M187 320 38 240 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=46900 $D=1
M188 6 319 729 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=42270 $D=1
M189 6 320 730 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=46900 $D=1
M190 321 729 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=42270 $D=1
M191 322 730 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=46900 $D=1
M192 319 315 321 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=42270 $D=1
M193 320 316 322 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=46900 $D=1
M194 321 39 249 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=42270 $D=1
M195 322 39 250 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=46900 $D=1
M196 253 40 321 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=42270 $D=1
M197 254 40 322 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=46900 $D=1
M198 323 40 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=42270 $D=1
M199 324 40 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=46900 $D=1
M200 6 41 325 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=42270 $D=1
M201 6 41 326 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=46900 $D=1
M202 327 42 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=42270 $D=1
M203 328 42 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=46900 $D=1
M204 329 41 239 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=42270 $D=1
M205 330 41 240 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=46900 $D=1
M206 6 329 731 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=42270 $D=1
M207 6 330 732 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=46900 $D=1
M208 331 731 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=42270 $D=1
M209 332 732 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=46900 $D=1
M210 329 325 331 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=42270 $D=1
M211 330 326 332 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=46900 $D=1
M212 331 42 249 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=42270 $D=1
M213 332 42 250 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=46900 $D=1
M214 253 43 331 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=42270 $D=1
M215 254 43 332 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=46900 $D=1
M216 333 43 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=42270 $D=1
M217 334 43 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=46900 $D=1
M218 6 44 335 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=42270 $D=1
M219 6 44 336 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=46900 $D=1
M220 337 45 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=42270 $D=1
M221 338 45 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=46900 $D=1
M222 339 44 239 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=42270 $D=1
M223 340 44 240 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=46900 $D=1
M224 6 339 733 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=42270 $D=1
M225 6 340 734 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=46900 $D=1
M226 341 733 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=42270 $D=1
M227 342 734 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=46900 $D=1
M228 339 335 341 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=42270 $D=1
M229 340 336 342 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=46900 $D=1
M230 341 45 249 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=42270 $D=1
M231 342 45 250 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=46900 $D=1
M232 253 46 341 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=42270 $D=1
M233 254 46 342 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=46900 $D=1
M234 343 46 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=42270 $D=1
M235 344 46 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=46900 $D=1
M236 6 47 345 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=42270 $D=1
M237 6 47 346 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=46900 $D=1
M238 347 48 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=42270 $D=1
M239 348 48 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=46900 $D=1
M240 349 47 239 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=42270 $D=1
M241 350 47 240 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=46900 $D=1
M242 6 349 735 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=42270 $D=1
M243 6 350 736 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=46900 $D=1
M244 351 735 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=42270 $D=1
M245 352 736 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=46900 $D=1
M246 349 345 351 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=42270 $D=1
M247 350 346 352 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=46900 $D=1
M248 351 48 249 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=42270 $D=1
M249 352 48 250 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=46900 $D=1
M250 253 49 351 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=42270 $D=1
M251 254 49 352 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=46900 $D=1
M252 353 49 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=42270 $D=1
M253 354 49 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=46900 $D=1
M254 6 50 355 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=42270 $D=1
M255 6 50 356 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=46900 $D=1
M256 357 51 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=42270 $D=1
M257 358 51 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=46900 $D=1
M258 359 50 239 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=42270 $D=1
M259 360 50 240 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=46900 $D=1
M260 6 359 737 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=42270 $D=1
M261 6 360 738 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=46900 $D=1
M262 361 737 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=42270 $D=1
M263 362 738 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=46900 $D=1
M264 359 355 361 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=42270 $D=1
M265 360 356 362 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=46900 $D=1
M266 361 51 249 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=42270 $D=1
M267 362 51 250 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=46900 $D=1
M268 253 52 361 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=42270 $D=1
M269 254 52 362 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=46900 $D=1
M270 363 52 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=42270 $D=1
M271 364 52 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=46900 $D=1
M272 6 53 365 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=42270 $D=1
M273 6 53 366 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=46900 $D=1
M274 367 54 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=42270 $D=1
M275 368 54 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=46900 $D=1
M276 369 53 239 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=42270 $D=1
M277 370 53 240 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=46900 $D=1
M278 6 369 739 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=42270 $D=1
M279 6 370 740 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=46900 $D=1
M280 371 739 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=42270 $D=1
M281 372 740 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=46900 $D=1
M282 369 365 371 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=42270 $D=1
M283 370 366 372 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=46900 $D=1
M284 371 54 249 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=42270 $D=1
M285 372 54 250 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=46900 $D=1
M286 253 55 371 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=42270 $D=1
M287 254 55 372 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=46900 $D=1
M288 373 55 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=42270 $D=1
M289 374 55 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=46900 $D=1
M290 6 56 375 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=42270 $D=1
M291 6 56 376 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=46900 $D=1
M292 377 57 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=42270 $D=1
M293 378 57 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=46900 $D=1
M294 379 56 239 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=42270 $D=1
M295 380 56 240 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=46900 $D=1
M296 6 379 741 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=42270 $D=1
M297 6 380 742 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=46900 $D=1
M298 381 741 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=42270 $D=1
M299 382 742 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=46900 $D=1
M300 379 375 381 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=42270 $D=1
M301 380 376 382 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=46900 $D=1
M302 381 57 249 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=42270 $D=1
M303 382 57 250 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=46900 $D=1
M304 253 58 381 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=42270 $D=1
M305 254 58 382 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=46900 $D=1
M306 383 58 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=42270 $D=1
M307 384 58 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=46900 $D=1
M308 6 59 385 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=42270 $D=1
M309 6 59 386 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=46900 $D=1
M310 387 60 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=42270 $D=1
M311 388 60 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=46900 $D=1
M312 389 59 239 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=42270 $D=1
M313 390 59 240 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=46900 $D=1
M314 6 389 743 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=42270 $D=1
M315 6 390 744 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=46900 $D=1
M316 391 743 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=42270 $D=1
M317 392 744 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=46900 $D=1
M318 389 385 391 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=42270 $D=1
M319 390 386 392 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=46900 $D=1
M320 391 60 249 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=42270 $D=1
M321 392 60 250 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=46900 $D=1
M322 253 61 391 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=42270 $D=1
M323 254 61 392 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=46900 $D=1
M324 393 61 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=42270 $D=1
M325 394 61 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=46900 $D=1
M326 6 62 395 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=42270 $D=1
M327 6 62 396 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=46900 $D=1
M328 397 63 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=42270 $D=1
M329 398 63 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=46900 $D=1
M330 399 62 239 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=42270 $D=1
M331 400 62 240 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=46900 $D=1
M332 6 399 745 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=42270 $D=1
M333 6 400 746 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=46900 $D=1
M334 401 745 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=42270 $D=1
M335 402 746 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=46900 $D=1
M336 399 395 401 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=42270 $D=1
M337 400 396 402 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=46900 $D=1
M338 401 63 249 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=42270 $D=1
M339 402 63 250 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=46900 $D=1
M340 253 64 401 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=42270 $D=1
M341 254 64 402 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=46900 $D=1
M342 403 64 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=42270 $D=1
M343 404 64 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=46900 $D=1
M344 6 65 405 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=42270 $D=1
M345 6 65 406 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=46900 $D=1
M346 407 66 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=42270 $D=1
M347 408 66 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=46900 $D=1
M348 409 65 239 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=42270 $D=1
M349 410 65 240 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=46900 $D=1
M350 6 409 747 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=42270 $D=1
M351 6 410 748 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=46900 $D=1
M352 411 747 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=42270 $D=1
M353 412 748 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=46900 $D=1
M354 409 405 411 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=42270 $D=1
M355 410 406 412 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=46900 $D=1
M356 411 66 249 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=42270 $D=1
M357 412 66 250 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=46900 $D=1
M358 253 67 411 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=42270 $D=1
M359 254 67 412 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=46900 $D=1
M360 413 67 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=42270 $D=1
M361 414 67 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=46900 $D=1
M362 6 68 415 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=42270 $D=1
M363 6 68 416 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=46900 $D=1
M364 417 69 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=42270 $D=1
M365 418 69 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=46900 $D=1
M366 419 68 239 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=42270 $D=1
M367 420 68 240 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=46900 $D=1
M368 6 419 749 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=42270 $D=1
M369 6 420 750 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=46900 $D=1
M370 421 749 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=42270 $D=1
M371 422 750 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=46900 $D=1
M372 419 415 421 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=42270 $D=1
M373 420 416 422 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=46900 $D=1
M374 421 69 249 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=42270 $D=1
M375 422 69 250 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=46900 $D=1
M376 253 70 421 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=42270 $D=1
M377 254 70 422 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=46900 $D=1
M378 423 70 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=42270 $D=1
M379 424 70 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=46900 $D=1
M380 6 71 425 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=42270 $D=1
M381 6 71 426 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=46900 $D=1
M382 427 72 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=42270 $D=1
M383 428 72 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=46900 $D=1
M384 429 71 239 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=42270 $D=1
M385 430 71 240 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=46900 $D=1
M386 6 429 751 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=42270 $D=1
M387 6 430 752 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=46900 $D=1
M388 431 751 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=42270 $D=1
M389 432 752 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=46900 $D=1
M390 429 425 431 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=42270 $D=1
M391 430 426 432 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=46900 $D=1
M392 431 72 249 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=42270 $D=1
M393 432 72 250 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=46900 $D=1
M394 253 73 431 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=42270 $D=1
M395 254 73 432 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=46900 $D=1
M396 433 73 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=42270 $D=1
M397 434 73 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=46900 $D=1
M398 6 74 435 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=42270 $D=1
M399 6 74 436 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=46900 $D=1
M400 437 75 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=42270 $D=1
M401 438 75 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=46900 $D=1
M402 439 74 239 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=42270 $D=1
M403 440 74 240 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=46900 $D=1
M404 6 439 753 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=42270 $D=1
M405 6 440 754 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=46900 $D=1
M406 441 753 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=42270 $D=1
M407 442 754 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=46900 $D=1
M408 439 435 441 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=42270 $D=1
M409 440 436 442 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=46900 $D=1
M410 441 75 249 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=42270 $D=1
M411 442 75 250 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=46900 $D=1
M412 253 76 441 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=42270 $D=1
M413 254 76 442 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=46900 $D=1
M414 443 76 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=42270 $D=1
M415 444 76 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=46900 $D=1
M416 6 77 445 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=42270 $D=1
M417 6 77 446 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=46900 $D=1
M418 447 78 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=42270 $D=1
M419 448 78 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=46900 $D=1
M420 449 77 239 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=42270 $D=1
M421 450 77 240 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=46900 $D=1
M422 6 449 755 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=42270 $D=1
M423 6 450 756 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=46900 $D=1
M424 451 755 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=42270 $D=1
M425 452 756 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=46900 $D=1
M426 449 445 451 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=42270 $D=1
M427 450 446 452 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=46900 $D=1
M428 451 78 249 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=42270 $D=1
M429 452 78 250 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=46900 $D=1
M430 253 79 451 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=42270 $D=1
M431 254 79 452 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=46900 $D=1
M432 453 79 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=42270 $D=1
M433 454 79 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=46900 $D=1
M434 6 80 455 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=42270 $D=1
M435 6 80 456 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=46900 $D=1
M436 457 81 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=42270 $D=1
M437 458 81 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=46900 $D=1
M438 459 80 239 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=42270 $D=1
M439 460 80 240 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=46900 $D=1
M440 6 459 757 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=42270 $D=1
M441 6 460 758 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=46900 $D=1
M442 461 757 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=42270 $D=1
M443 462 758 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=46900 $D=1
M444 459 455 461 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=42270 $D=1
M445 460 456 462 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=46900 $D=1
M446 461 81 249 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=42270 $D=1
M447 462 81 250 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=46900 $D=1
M448 253 82 461 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=42270 $D=1
M449 254 82 462 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=46900 $D=1
M450 463 82 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=42270 $D=1
M451 464 82 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=46900 $D=1
M452 6 83 465 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=42270 $D=1
M453 6 83 466 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=46900 $D=1
M454 467 84 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=42270 $D=1
M455 468 84 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=46900 $D=1
M456 469 83 239 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=42270 $D=1
M457 470 83 240 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=46900 $D=1
M458 6 469 759 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=42270 $D=1
M459 6 470 760 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=46900 $D=1
M460 471 759 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=42270 $D=1
M461 472 760 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=46900 $D=1
M462 469 465 471 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=42270 $D=1
M463 470 466 472 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=46900 $D=1
M464 471 84 249 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=42270 $D=1
M465 472 84 250 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=46900 $D=1
M466 253 85 471 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=42270 $D=1
M467 254 85 472 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=46900 $D=1
M468 473 85 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=42270 $D=1
M469 474 85 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=46900 $D=1
M470 6 86 475 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=42270 $D=1
M471 6 86 476 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=46900 $D=1
M472 477 87 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=42270 $D=1
M473 478 87 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=46900 $D=1
M474 479 86 239 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=42270 $D=1
M475 480 86 240 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=46900 $D=1
M476 6 479 761 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=42270 $D=1
M477 6 480 762 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=46900 $D=1
M478 481 761 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=42270 $D=1
M479 482 762 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=46900 $D=1
M480 479 475 481 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=42270 $D=1
M481 480 476 482 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=46900 $D=1
M482 481 87 249 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=42270 $D=1
M483 482 87 250 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=46900 $D=1
M484 253 88 481 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=42270 $D=1
M485 254 88 482 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=46900 $D=1
M486 483 88 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=42270 $D=1
M487 484 88 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=46900 $D=1
M488 6 89 485 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=42270 $D=1
M489 6 89 486 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=46900 $D=1
M490 487 90 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=42270 $D=1
M491 488 90 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=46900 $D=1
M492 489 89 239 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=42270 $D=1
M493 490 89 240 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=46900 $D=1
M494 6 489 763 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=42270 $D=1
M495 6 490 764 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=46900 $D=1
M496 491 763 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=42270 $D=1
M497 492 764 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=46900 $D=1
M498 489 485 491 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=42270 $D=1
M499 490 486 492 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=46900 $D=1
M500 491 90 249 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=42270 $D=1
M501 492 90 250 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=46900 $D=1
M502 253 91 491 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=42270 $D=1
M503 254 91 492 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=46900 $D=1
M504 493 91 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=42270 $D=1
M505 494 91 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=46900 $D=1
M506 6 92 495 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=42270 $D=1
M507 6 92 496 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=46900 $D=1
M508 497 93 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=42270 $D=1
M509 498 93 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=46900 $D=1
M510 499 92 239 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=42270 $D=1
M511 500 92 240 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=46900 $D=1
M512 6 499 765 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=42270 $D=1
M513 6 500 766 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=46900 $D=1
M514 501 765 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=42270 $D=1
M515 502 766 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=46900 $D=1
M516 499 495 501 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=42270 $D=1
M517 500 496 502 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=46900 $D=1
M518 501 93 249 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=42270 $D=1
M519 502 93 250 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=46900 $D=1
M520 253 94 501 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=42270 $D=1
M521 254 94 502 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=46900 $D=1
M522 503 94 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=42270 $D=1
M523 504 94 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=46900 $D=1
M524 6 95 505 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=42270 $D=1
M525 6 95 506 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=46900 $D=1
M526 507 96 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=42270 $D=1
M527 508 96 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=46900 $D=1
M528 509 95 239 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=42270 $D=1
M529 510 95 240 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=46900 $D=1
M530 6 509 767 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=42270 $D=1
M531 6 510 768 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=46900 $D=1
M532 511 767 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=42270 $D=1
M533 512 768 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=46900 $D=1
M534 509 505 511 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=42270 $D=1
M535 510 506 512 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=46900 $D=1
M536 511 96 249 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=42270 $D=1
M537 512 96 250 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=46900 $D=1
M538 253 97 511 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=42270 $D=1
M539 254 97 512 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=46900 $D=1
M540 513 97 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=42270 $D=1
M541 514 97 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=46900 $D=1
M542 6 98 515 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=42270 $D=1
M543 6 98 516 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=46900 $D=1
M544 517 99 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=42270 $D=1
M545 518 99 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=46900 $D=1
M546 519 98 239 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=42270 $D=1
M547 520 98 240 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=46900 $D=1
M548 6 519 769 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=42270 $D=1
M549 6 520 770 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=46900 $D=1
M550 521 769 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=42270 $D=1
M551 522 770 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=46900 $D=1
M552 519 515 521 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=42270 $D=1
M553 520 516 522 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=46900 $D=1
M554 521 99 249 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=42270 $D=1
M555 522 99 250 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=46900 $D=1
M556 253 100 521 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=42270 $D=1
M557 254 100 522 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=46900 $D=1
M558 523 100 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=42270 $D=1
M559 524 100 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=46900 $D=1
M560 6 101 525 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=42270 $D=1
M561 6 101 526 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=46900 $D=1
M562 527 102 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=42270 $D=1
M563 528 102 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=46900 $D=1
M564 529 101 239 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=42270 $D=1
M565 530 101 240 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=46900 $D=1
M566 6 529 771 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=42270 $D=1
M567 6 530 772 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=46900 $D=1
M568 531 771 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=42270 $D=1
M569 532 772 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=46900 $D=1
M570 529 525 531 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=42270 $D=1
M571 530 526 532 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=46900 $D=1
M572 531 102 249 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=42270 $D=1
M573 532 102 250 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=46900 $D=1
M574 253 103 531 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=42270 $D=1
M575 254 103 532 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=46900 $D=1
M576 533 103 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=42270 $D=1
M577 534 103 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=46900 $D=1
M578 6 104 535 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=42270 $D=1
M579 6 104 536 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=46900 $D=1
M580 537 105 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=42270 $D=1
M581 538 105 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=46900 $D=1
M582 539 104 239 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=42270 $D=1
M583 540 104 240 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=46900 $D=1
M584 6 539 773 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=42270 $D=1
M585 6 540 774 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=46900 $D=1
M586 541 773 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=42270 $D=1
M587 542 774 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=46900 $D=1
M588 539 535 541 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=42270 $D=1
M589 540 536 542 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=46900 $D=1
M590 541 105 249 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=42270 $D=1
M591 542 105 250 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=46900 $D=1
M592 253 109 541 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=42270 $D=1
M593 254 109 542 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=46900 $D=1
M594 543 109 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=42270 $D=1
M595 544 109 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=46900 $D=1
M596 6 110 545 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=42270 $D=1
M597 6 110 546 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=46900 $D=1
M598 547 111 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=42270 $D=1
M599 548 111 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=46900 $D=1
M600 549 110 239 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=42270 $D=1
M601 550 110 240 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=46900 $D=1
M602 6 549 775 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=42270 $D=1
M603 6 550 776 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=46900 $D=1
M604 551 775 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=42270 $D=1
M605 552 776 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=46900 $D=1
M606 549 545 551 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=42270 $D=1
M607 550 546 552 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=46900 $D=1
M608 551 111 249 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=42270 $D=1
M609 552 111 250 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=46900 $D=1
M610 253 113 551 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=42270 $D=1
M611 254 113 552 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=46900 $D=1
M612 553 113 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=42270 $D=1
M613 554 113 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=46900 $D=1
M614 6 114 555 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=42270 $D=1
M615 6 114 556 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=46900 $D=1
M616 557 115 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=42270 $D=1
M617 558 115 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=46900 $D=1
M618 6 115 249 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=42270 $D=1
M619 6 115 250 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=46900 $D=1
M620 253 114 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=42270 $D=1
M621 254 114 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=46900 $D=1
M622 6 561 559 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=42270 $D=1
M623 6 562 560 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=46900 $D=1
M624 561 117 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=42270 $D=1
M625 562 117 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=46900 $D=1
M626 777 249 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=42270 $D=1
M627 778 250 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=46900 $D=1
M628 563 559 777 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=42270 $D=1
M629 564 560 778 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=46900 $D=1
M630 6 563 565 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=42270 $D=1
M631 6 564 566 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=46900 $D=1
M632 779 565 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=42270 $D=1
M633 780 566 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=46900 $D=1
M634 563 561 779 6 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=42270 $D=1
M635 564 562 780 6 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=46900 $D=1
M636 6 569 567 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=42270 $D=1
M637 6 570 568 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=46900 $D=1
M638 569 117 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=42270 $D=1
M639 570 117 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=46900 $D=1
M640 781 253 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=42270 $D=1
M641 782 254 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=46900 $D=1
M642 571 567 781 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=42270 $D=1
M643 572 568 782 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=46900 $D=1
M644 6 571 119 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=42270 $D=1
M645 6 572 120 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=46900 $D=1
M646 783 119 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=42270 $D=1
M647 784 120 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=46900 $D=1
M648 571 569 783 6 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=42270 $D=1
M649 572 570 784 6 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=46900 $D=1
M650 573 121 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=42270 $D=1
M651 574 121 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=46900 $D=1
M652 575 573 565 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=42270 $D=1
M653 576 574 566 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=46900 $D=1
M654 122 121 575 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=42270 $D=1
M655 123 121 576 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=46900 $D=1
M656 577 124 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=42270 $D=1
M657 578 124 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=46900 $D=1
M658 579 577 119 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=42270 $D=1
M659 580 578 120 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=46900 $D=1
M660 785 124 579 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=42270 $D=1
M661 786 124 580 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=46900 $D=1
M662 6 119 785 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=42270 $D=1
M663 6 120 786 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=46900 $D=1
M664 581 125 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=42270 $D=1
M665 582 125 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=46900 $D=1
M666 583 581 579 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=42270 $D=1
M667 584 582 580 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=46900 $D=1
M668 11 125 583 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=42270 $D=1
M669 12 125 584 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=46900 $D=1
M670 586 585 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=42270 $D=1
M671 587 126 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=46900 $D=1
M672 6 590 588 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=42270 $D=1
M673 6 591 589 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=46900 $D=1
M674 592 575 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=42270 $D=1
M675 593 576 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=46900 $D=1
M676 590 592 585 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=42270 $D=1
M677 591 593 126 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=46900 $D=1
M678 586 575 590 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=42270 $D=1
M679 587 576 591 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=46900 $D=1
M680 594 588 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=42270 $D=1
M681 595 589 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=46900 $D=1
M682 127 594 583 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=42270 $D=1
M683 585 595 584 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=46900 $D=1
M684 575 588 127 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=42270 $D=1
M685 576 589 585 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=46900 $D=1
M686 596 127 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=42270 $D=1
M687 597 585 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=46900 $D=1
M688 598 588 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=42270 $D=1
M689 599 589 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=46900 $D=1
M690 600 598 596 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=42270 $D=1
M691 601 599 597 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=46900 $D=1
M692 583 588 600 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=42270 $D=1
M693 584 589 601 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=46900 $D=1
M694 602 575 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=42270 $D=1
M695 603 576 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=46900 $D=1
M696 6 583 602 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=42270 $D=1
M697 6 584 603 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=46900 $D=1
M698 604 600 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=42270 $D=1
M699 605 601 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=46900 $D=1
M700 805 575 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=42270 $D=1
M701 806 576 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=46900 $D=1
M702 606 583 805 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=42270 $D=1
M703 607 584 806 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=46900 $D=1
M704 807 575 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=42270 $D=1
M705 808 576 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=46900 $D=1
M706 608 583 807 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=42270 $D=1
M707 609 584 808 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=46900 $D=1
M708 612 575 610 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=42270 $D=1
M709 613 576 611 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=46900 $D=1
M710 610 583 612 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=42270 $D=1
M711 611 584 613 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=46900 $D=1
M712 6 608 610 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=42270 $D=1
M713 6 609 611 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=46900 $D=1
M714 614 130 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=42270 $D=1
M715 615 130 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=46900 $D=1
M716 616 614 602 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=42270 $D=1
M717 617 615 603 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=46900 $D=1
M718 606 130 616 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=42270 $D=1
M719 607 130 617 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=46900 $D=1
M720 618 614 604 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=42270 $D=1
M721 619 615 605 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=46900 $D=1
M722 612 130 618 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=42270 $D=1
M723 613 130 619 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=46900 $D=1
M724 620 131 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=42270 $D=1
M725 621 131 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=46900 $D=1
M726 622 620 618 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=42270 $D=1
M727 623 621 619 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=46900 $D=1
M728 616 131 622 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=42270 $D=1
M729 617 131 623 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=46900 $D=1
M730 13 622 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=42270 $D=1
M731 14 623 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=46900 $D=1
M732 624 132 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=42270 $D=1
M733 625 132 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=46900 $D=1
M734 626 624 133 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=42270 $D=1
M735 627 625 134 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=46900 $D=1
M736 135 132 626 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=42270 $D=1
M737 136 132 627 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=46900 $D=1
M738 628 132 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=42270 $D=1
M739 629 132 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=46900 $D=1
M740 630 628 137 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=42270 $D=1
M741 631 629 138 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=46900 $D=1
M742 139 132 630 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=42270 $D=1
M743 140 132 631 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=46900 $D=1
M744 632 132 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=42270 $D=1
M745 633 132 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=46900 $D=1
M746 634 632 129 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=42270 $D=1
M747 635 633 128 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=46900 $D=1
M748 141 132 634 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=42270 $D=1
M749 108 132 635 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=46900 $D=1
M750 636 132 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=42270 $D=1
M751 637 132 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=46900 $D=1
M752 638 636 142 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=42270 $D=1
M753 639 637 143 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=46900 $D=1
M754 144 132 638 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=42270 $D=1
M755 145 132 639 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=46900 $D=1
M756 640 132 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=42270 $D=1
M757 641 132 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=46900 $D=1
M758 642 640 146 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=42270 $D=1
M759 643 641 147 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=46900 $D=1
M760 148 132 642 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=42270 $D=1
M761 148 132 643 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=46900 $D=1
M762 6 575 787 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=42270 $D=1
M763 6 576 788 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=46900 $D=1
M764 136 787 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=42270 $D=1
M765 133 788 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=46900 $D=1
M766 644 149 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=42270 $D=1
M767 645 149 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=46900 $D=1
M768 150 644 136 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=42270 $D=1
M769 151 645 133 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=46900 $D=1
M770 626 149 150 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=42270 $D=1
M771 627 149 151 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=46900 $D=1
M772 646 152 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=42270 $D=1
M773 647 152 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=46900 $D=1
M774 153 646 150 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=42270 $D=1
M775 116 647 151 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=46900 $D=1
M776 630 152 153 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=42270 $D=1
M777 631 152 116 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=46900 $D=1
M778 648 154 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=42270 $D=1
M779 649 154 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=46900 $D=1
M780 155 648 153 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=42270 $D=1
M781 106 649 116 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=46900 $D=1
M782 634 154 155 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=42270 $D=1
M783 635 154 106 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=46900 $D=1
M784 650 156 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=42270 $D=1
M785 651 156 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=46900 $D=1
M786 157 650 155 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=42270 $D=1
M787 158 651 106 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=46900 $D=1
M788 638 156 157 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=42270 $D=1
M789 639 156 158 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=46900 $D=1
M790 652 159 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=42270 $D=1
M791 653 159 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=46900 $D=1
M792 225 652 157 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=42270 $D=1
M793 226 653 158 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=46900 $D=1
M794 642 159 225 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=42270 $D=1
M795 643 159 226 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=46900 $D=1
M796 654 160 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=42270 $D=1
M797 655 160 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=46900 $D=1
M798 656 654 119 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=42270 $D=1
M799 657 655 120 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=46900 $D=1
M800 11 160 656 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=42270 $D=1
M801 12 160 657 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=46900 $D=1
M802 809 565 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=42270 $D=1
M803 810 566 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=46900 $D=1
M804 658 656 809 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=42270 $D=1
M805 659 657 810 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=46900 $D=1
M806 662 565 660 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=42270 $D=1
M807 663 566 661 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=46900 $D=1
M808 660 656 662 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=42270 $D=1
M809 661 657 663 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=46900 $D=1
M810 6 658 660 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=42270 $D=1
M811 6 659 661 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=46900 $D=1
M812 811 161 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=42270 $D=1
M813 812 664 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=46900 $D=1
M814 789 662 811 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=42270 $D=1
M815 790 663 812 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=46900 $D=1
M816 664 789 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=42270 $D=1
M817 162 790 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=46900 $D=1
M818 665 565 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=42270 $D=1
M819 666 566 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=46900 $D=1
M820 6 667 665 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=42270 $D=1
M821 6 668 666 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=46900 $D=1
M822 667 656 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=42270 $D=1
M823 668 657 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=46900 $D=1
M824 813 665 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=42270 $D=1
M825 814 666 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=46900 $D=1
M826 669 161 813 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=42270 $D=1
M827 670 664 814 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=46900 $D=1
M828 672 163 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=42270 $D=1
M829 673 671 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=46900 $D=1
M830 815 669 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=42270 $D=1
M831 816 670 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=46900 $D=1
M832 671 672 815 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=42270 $D=1
M833 164 673 816 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=46900 $D=1
M834 675 674 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=42270 $D=1
M835 676 165 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=46900 $D=1
M836 6 679 677 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=42270 $D=1
M837 6 680 678 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=46900 $D=1
M838 681 122 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=42270 $D=1
M839 682 123 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=46900 $D=1
M840 679 681 674 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=42270 $D=1
M841 680 682 165 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=46900 $D=1
M842 675 122 679 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=42270 $D=1
M843 676 123 680 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=46900 $D=1
M844 683 677 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=42270 $D=1
M845 684 678 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=46900 $D=1
M846 166 683 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=42270 $D=1
M847 674 684 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=46900 $D=1
M848 122 677 166 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=42270 $D=1
M849 123 678 674 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=46900 $D=1
M850 685 166 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=42270 $D=1
M851 686 674 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=46900 $D=1
M852 687 677 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=42270 $D=1
M853 688 678 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=46900 $D=1
M854 227 687 685 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=42270 $D=1
M855 228 688 686 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=46900 $D=1
M856 6 677 227 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=42270 $D=1
M857 6 678 228 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=46900 $D=1
M858 689 167 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=42270 $D=1
M859 690 167 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=46900 $D=1
M860 691 689 227 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=42270 $D=1
M861 692 690 228 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=46900 $D=1
M862 13 167 691 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=42270 $D=1
M863 14 167 692 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=46900 $D=1
M864 693 168 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=42270 $D=1
M865 694 168 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=46900 $D=1
M866 695 693 691 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=42270 $D=1
M867 696 694 692 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=46900 $D=1
M868 6 168 695 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=42270 $D=1
M869 6 168 696 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=46900 $D=1
M870 697 117 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=42270 $D=1
M871 698 117 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=46900 $D=1
M872 6 697 699 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=42270 $D=1
M873 6 698 700 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=46900 $D=1
M874 701 117 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=42270 $D=1
M875 702 117 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=46900 $D=1
M876 703 697 695 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=42270 $D=1
M877 704 698 696 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=46900 $D=1
M878 6 703 791 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=42270 $D=1
M879 6 704 792 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=46900 $D=1
M880 705 791 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=42270 $D=1
M881 706 792 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=46900 $D=1
M882 703 699 705 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=42270 $D=1
M883 704 700 706 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=46900 $D=1
M884 707 117 705 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=42270 $D=1
M885 708 117 706 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=46900 $D=1
M886 6 711 709 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=42270 $D=1
M887 6 712 710 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=46900 $D=1
M888 711 117 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=42270 $D=1
M889 712 117 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=46900 $D=1
M890 793 707 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=42270 $D=1
M891 794 708 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=46900 $D=1
M892 713 709 793 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=42270 $D=1
M893 714 710 794 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=46900 $D=1
M894 6 713 122 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=42270 $D=1
M895 6 714 123 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=46900 $D=1
M896 795 122 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=42270 $D=1
M897 796 123 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=46900 $D=1
M898 713 711 795 6 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=42270 $D=1
M899 714 712 796 6 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=46900 $D=1
M900 201 1 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=43520 $D=0
M901 202 1 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=48150 $D=0
M902 203 1 2 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=43520 $D=0
M903 204 1 3 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=48150 $D=0
M904 6 201 203 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=43520 $D=0
M905 6 202 204 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=48150 $D=0
M906 205 1 4 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=43520 $D=0
M907 206 1 4 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=48150 $D=0
M908 5 201 205 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=43520 $D=0
M909 5 202 206 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=48150 $D=0
M910 207 1 6 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=43520 $D=0
M911 208 1 6 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=48150 $D=0
M912 6 201 207 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=43520 $D=0
M913 6 202 208 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=48150 $D=0
M914 211 7 207 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=43520 $D=0
M915 212 7 208 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=48150 $D=0
M916 209 7 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=43520 $D=0
M917 210 7 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=48150 $D=0
M918 213 7 205 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=43520 $D=0
M919 214 7 206 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=48150 $D=0
M920 203 209 213 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=43520 $D=0
M921 204 210 214 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=48150 $D=0
M922 215 8 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=43520 $D=0
M923 216 8 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=48150 $D=0
M924 217 8 213 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=43520 $D=0
M925 218 8 214 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=48150 $D=0
M926 211 215 217 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=43520 $D=0
M927 212 216 218 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=48150 $D=0
M928 219 10 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=43520 $D=0
M929 220 10 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=48150 $D=0
M930 221 10 6 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=43520 $D=0
M931 222 10 6 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=48150 $D=0
M932 11 219 221 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=43520 $D=0
M933 12 220 222 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=48150 $D=0
M934 223 10 13 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=43520 $D=0
M935 224 10 14 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=48150 $D=0
M936 225 219 223 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=43520 $D=0
M937 226 220 224 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=48150 $D=0
M938 229 10 227 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=43520 $D=0
M939 230 10 228 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=48150 $D=0
M940 217 219 229 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=43520 $D=0
M941 218 220 230 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=48150 $D=0
M942 233 15 229 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=43520 $D=0
M943 234 15 230 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=48150 $D=0
M944 231 15 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=43520 $D=0
M945 232 15 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=48150 $D=0
M946 235 15 223 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=43520 $D=0
M947 236 15 224 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=48150 $D=0
M948 221 231 235 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=43520 $D=0
M949 222 232 236 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=48150 $D=0
M950 237 16 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=43520 $D=0
M951 238 16 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=48150 $D=0
M952 239 16 235 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=43520 $D=0
M953 240 16 236 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=48150 $D=0
M954 233 237 239 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=43520 $D=0
M955 234 238 240 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=48150 $D=0
M956 9 17 241 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=43520 $D=0
M957 9 17 242 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=48150 $D=0
M958 243 18 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=43520 $D=0
M959 244 18 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=48150 $D=0
M960 245 241 239 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=43520 $D=0
M961 246 242 240 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=48150 $D=0
M962 9 245 715 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=43520 $D=0
M963 9 246 716 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=48150 $D=0
M964 247 715 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=43520 $D=0
M965 248 716 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=48150 $D=0
M966 245 17 247 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=43520 $D=0
M967 246 17 248 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=48150 $D=0
M968 247 243 249 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=43520 $D=0
M969 248 244 250 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=48150 $D=0
M970 253 251 247 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=43520 $D=0
M971 254 252 248 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=48150 $D=0
M972 251 19 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=43520 $D=0
M973 252 19 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=48150 $D=0
M974 9 20 255 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=43520 $D=0
M975 9 20 256 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=48150 $D=0
M976 257 21 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=43520 $D=0
M977 258 21 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=48150 $D=0
M978 259 255 239 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=43520 $D=0
M979 260 256 240 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=48150 $D=0
M980 9 259 717 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=43520 $D=0
M981 9 260 718 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=48150 $D=0
M982 261 717 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=43520 $D=0
M983 262 718 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=48150 $D=0
M984 259 20 261 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=43520 $D=0
M985 260 20 262 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=48150 $D=0
M986 261 257 249 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=43520 $D=0
M987 262 258 250 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=48150 $D=0
M988 253 263 261 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=43520 $D=0
M989 254 264 262 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=48150 $D=0
M990 263 22 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=43520 $D=0
M991 264 22 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=48150 $D=0
M992 9 23 265 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=43520 $D=0
M993 9 23 266 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=48150 $D=0
M994 267 24 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=43520 $D=0
M995 268 24 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=48150 $D=0
M996 269 265 239 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=43520 $D=0
M997 270 266 240 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=48150 $D=0
M998 9 269 719 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=43520 $D=0
M999 9 270 720 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=48150 $D=0
M1000 271 719 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=43520 $D=0
M1001 272 720 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=48150 $D=0
M1002 269 23 271 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=43520 $D=0
M1003 270 23 272 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=48150 $D=0
M1004 271 267 249 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=43520 $D=0
M1005 272 268 250 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=48150 $D=0
M1006 253 273 271 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=43520 $D=0
M1007 254 274 272 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=48150 $D=0
M1008 273 25 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=43520 $D=0
M1009 274 25 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=48150 $D=0
M1010 9 26 275 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=43520 $D=0
M1011 9 26 276 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=48150 $D=0
M1012 277 27 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=43520 $D=0
M1013 278 27 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=48150 $D=0
M1014 279 275 239 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=43520 $D=0
M1015 280 276 240 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=48150 $D=0
M1016 9 279 721 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=43520 $D=0
M1017 9 280 722 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=48150 $D=0
M1018 281 721 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=43520 $D=0
M1019 282 722 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=48150 $D=0
M1020 279 26 281 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=43520 $D=0
M1021 280 26 282 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=48150 $D=0
M1022 281 277 249 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=43520 $D=0
M1023 282 278 250 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=48150 $D=0
M1024 253 283 281 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=43520 $D=0
M1025 254 284 282 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=48150 $D=0
M1026 283 28 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=43520 $D=0
M1027 284 28 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=48150 $D=0
M1028 9 29 285 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=43520 $D=0
M1029 9 29 286 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=48150 $D=0
M1030 287 30 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=43520 $D=0
M1031 288 30 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=48150 $D=0
M1032 289 285 239 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=43520 $D=0
M1033 290 286 240 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=48150 $D=0
M1034 9 289 723 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=43520 $D=0
M1035 9 290 724 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=48150 $D=0
M1036 291 723 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=43520 $D=0
M1037 292 724 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=48150 $D=0
M1038 289 29 291 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=43520 $D=0
M1039 290 29 292 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=48150 $D=0
M1040 291 287 249 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=43520 $D=0
M1041 292 288 250 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=48150 $D=0
M1042 253 293 291 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=43520 $D=0
M1043 254 294 292 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=48150 $D=0
M1044 293 31 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=43520 $D=0
M1045 294 31 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=48150 $D=0
M1046 9 32 295 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=43520 $D=0
M1047 9 32 296 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=48150 $D=0
M1048 297 33 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=43520 $D=0
M1049 298 33 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=48150 $D=0
M1050 299 295 239 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=43520 $D=0
M1051 300 296 240 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=48150 $D=0
M1052 9 299 725 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=43520 $D=0
M1053 9 300 726 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=48150 $D=0
M1054 301 725 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=43520 $D=0
M1055 302 726 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=48150 $D=0
M1056 299 32 301 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=43520 $D=0
M1057 300 32 302 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=48150 $D=0
M1058 301 297 249 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=43520 $D=0
M1059 302 298 250 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=48150 $D=0
M1060 253 303 301 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=43520 $D=0
M1061 254 304 302 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=48150 $D=0
M1062 303 34 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=43520 $D=0
M1063 304 34 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=48150 $D=0
M1064 9 35 305 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=43520 $D=0
M1065 9 35 306 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=48150 $D=0
M1066 307 36 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=43520 $D=0
M1067 308 36 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=48150 $D=0
M1068 309 305 239 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=43520 $D=0
M1069 310 306 240 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=48150 $D=0
M1070 9 309 727 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=43520 $D=0
M1071 9 310 728 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=48150 $D=0
M1072 311 727 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=43520 $D=0
M1073 312 728 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=48150 $D=0
M1074 309 35 311 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=43520 $D=0
M1075 310 35 312 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=48150 $D=0
M1076 311 307 249 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=43520 $D=0
M1077 312 308 250 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=48150 $D=0
M1078 253 313 311 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=43520 $D=0
M1079 254 314 312 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=48150 $D=0
M1080 313 37 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=43520 $D=0
M1081 314 37 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=48150 $D=0
M1082 9 38 315 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=43520 $D=0
M1083 9 38 316 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=48150 $D=0
M1084 317 39 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=43520 $D=0
M1085 318 39 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=48150 $D=0
M1086 319 315 239 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=43520 $D=0
M1087 320 316 240 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=48150 $D=0
M1088 9 319 729 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=43520 $D=0
M1089 9 320 730 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=48150 $D=0
M1090 321 729 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=43520 $D=0
M1091 322 730 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=48150 $D=0
M1092 319 38 321 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=43520 $D=0
M1093 320 38 322 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=48150 $D=0
M1094 321 317 249 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=43520 $D=0
M1095 322 318 250 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=48150 $D=0
M1096 253 323 321 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=43520 $D=0
M1097 254 324 322 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=48150 $D=0
M1098 323 40 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=43520 $D=0
M1099 324 40 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=48150 $D=0
M1100 9 41 325 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=43520 $D=0
M1101 9 41 326 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=48150 $D=0
M1102 327 42 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=43520 $D=0
M1103 328 42 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=48150 $D=0
M1104 329 325 239 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=43520 $D=0
M1105 330 326 240 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=48150 $D=0
M1106 9 329 731 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=43520 $D=0
M1107 9 330 732 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=48150 $D=0
M1108 331 731 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=43520 $D=0
M1109 332 732 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=48150 $D=0
M1110 329 41 331 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=43520 $D=0
M1111 330 41 332 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=48150 $D=0
M1112 331 327 249 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=43520 $D=0
M1113 332 328 250 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=48150 $D=0
M1114 253 333 331 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=43520 $D=0
M1115 254 334 332 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=48150 $D=0
M1116 333 43 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=43520 $D=0
M1117 334 43 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=48150 $D=0
M1118 9 44 335 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=43520 $D=0
M1119 9 44 336 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=48150 $D=0
M1120 337 45 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=43520 $D=0
M1121 338 45 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=48150 $D=0
M1122 339 335 239 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=43520 $D=0
M1123 340 336 240 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=48150 $D=0
M1124 9 339 733 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=43520 $D=0
M1125 9 340 734 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=48150 $D=0
M1126 341 733 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=43520 $D=0
M1127 342 734 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=48150 $D=0
M1128 339 44 341 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=43520 $D=0
M1129 340 44 342 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=48150 $D=0
M1130 341 337 249 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=43520 $D=0
M1131 342 338 250 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=48150 $D=0
M1132 253 343 341 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=43520 $D=0
M1133 254 344 342 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=48150 $D=0
M1134 343 46 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=43520 $D=0
M1135 344 46 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=48150 $D=0
M1136 9 47 345 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=43520 $D=0
M1137 9 47 346 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=48150 $D=0
M1138 347 48 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=43520 $D=0
M1139 348 48 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=48150 $D=0
M1140 349 345 239 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=43520 $D=0
M1141 350 346 240 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=48150 $D=0
M1142 9 349 735 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=43520 $D=0
M1143 9 350 736 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=48150 $D=0
M1144 351 735 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=43520 $D=0
M1145 352 736 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=48150 $D=0
M1146 349 47 351 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=43520 $D=0
M1147 350 47 352 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=48150 $D=0
M1148 351 347 249 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=43520 $D=0
M1149 352 348 250 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=48150 $D=0
M1150 253 353 351 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=43520 $D=0
M1151 254 354 352 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=48150 $D=0
M1152 353 49 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=43520 $D=0
M1153 354 49 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=48150 $D=0
M1154 9 50 355 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=43520 $D=0
M1155 9 50 356 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=48150 $D=0
M1156 357 51 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=43520 $D=0
M1157 358 51 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=48150 $D=0
M1158 359 355 239 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=43520 $D=0
M1159 360 356 240 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=48150 $D=0
M1160 9 359 737 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=43520 $D=0
M1161 9 360 738 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=48150 $D=0
M1162 361 737 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=43520 $D=0
M1163 362 738 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=48150 $D=0
M1164 359 50 361 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=43520 $D=0
M1165 360 50 362 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=48150 $D=0
M1166 361 357 249 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=43520 $D=0
M1167 362 358 250 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=48150 $D=0
M1168 253 363 361 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=43520 $D=0
M1169 254 364 362 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=48150 $D=0
M1170 363 52 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=43520 $D=0
M1171 364 52 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=48150 $D=0
M1172 9 53 365 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=43520 $D=0
M1173 9 53 366 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=48150 $D=0
M1174 367 54 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=43520 $D=0
M1175 368 54 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=48150 $D=0
M1176 369 365 239 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=43520 $D=0
M1177 370 366 240 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=48150 $D=0
M1178 9 369 739 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=43520 $D=0
M1179 9 370 740 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=48150 $D=0
M1180 371 739 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=43520 $D=0
M1181 372 740 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=48150 $D=0
M1182 369 53 371 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=43520 $D=0
M1183 370 53 372 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=48150 $D=0
M1184 371 367 249 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=43520 $D=0
M1185 372 368 250 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=48150 $D=0
M1186 253 373 371 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=43520 $D=0
M1187 254 374 372 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=48150 $D=0
M1188 373 55 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=43520 $D=0
M1189 374 55 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=48150 $D=0
M1190 9 56 375 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=43520 $D=0
M1191 9 56 376 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=48150 $D=0
M1192 377 57 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=43520 $D=0
M1193 378 57 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=48150 $D=0
M1194 379 375 239 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=43520 $D=0
M1195 380 376 240 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=48150 $D=0
M1196 9 379 741 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=43520 $D=0
M1197 9 380 742 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=48150 $D=0
M1198 381 741 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=43520 $D=0
M1199 382 742 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=48150 $D=0
M1200 379 56 381 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=43520 $D=0
M1201 380 56 382 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=48150 $D=0
M1202 381 377 249 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=43520 $D=0
M1203 382 378 250 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=48150 $D=0
M1204 253 383 381 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=43520 $D=0
M1205 254 384 382 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=48150 $D=0
M1206 383 58 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=43520 $D=0
M1207 384 58 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=48150 $D=0
M1208 9 59 385 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=43520 $D=0
M1209 9 59 386 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=48150 $D=0
M1210 387 60 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=43520 $D=0
M1211 388 60 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=48150 $D=0
M1212 389 385 239 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=43520 $D=0
M1213 390 386 240 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=48150 $D=0
M1214 9 389 743 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=43520 $D=0
M1215 9 390 744 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=48150 $D=0
M1216 391 743 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=43520 $D=0
M1217 392 744 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=48150 $D=0
M1218 389 59 391 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=43520 $D=0
M1219 390 59 392 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=48150 $D=0
M1220 391 387 249 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=43520 $D=0
M1221 392 388 250 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=48150 $D=0
M1222 253 393 391 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=43520 $D=0
M1223 254 394 392 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=48150 $D=0
M1224 393 61 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=43520 $D=0
M1225 394 61 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=48150 $D=0
M1226 9 62 395 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=43520 $D=0
M1227 9 62 396 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=48150 $D=0
M1228 397 63 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=43520 $D=0
M1229 398 63 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=48150 $D=0
M1230 399 395 239 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=43520 $D=0
M1231 400 396 240 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=48150 $D=0
M1232 9 399 745 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=43520 $D=0
M1233 9 400 746 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=48150 $D=0
M1234 401 745 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=43520 $D=0
M1235 402 746 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=48150 $D=0
M1236 399 62 401 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=43520 $D=0
M1237 400 62 402 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=48150 $D=0
M1238 401 397 249 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=43520 $D=0
M1239 402 398 250 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=48150 $D=0
M1240 253 403 401 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=43520 $D=0
M1241 254 404 402 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=48150 $D=0
M1242 403 64 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=43520 $D=0
M1243 404 64 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=48150 $D=0
M1244 9 65 405 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=43520 $D=0
M1245 9 65 406 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=48150 $D=0
M1246 407 66 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=43520 $D=0
M1247 408 66 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=48150 $D=0
M1248 409 405 239 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=43520 $D=0
M1249 410 406 240 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=48150 $D=0
M1250 9 409 747 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=43520 $D=0
M1251 9 410 748 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=48150 $D=0
M1252 411 747 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=43520 $D=0
M1253 412 748 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=48150 $D=0
M1254 409 65 411 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=43520 $D=0
M1255 410 65 412 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=48150 $D=0
M1256 411 407 249 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=43520 $D=0
M1257 412 408 250 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=48150 $D=0
M1258 253 413 411 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=43520 $D=0
M1259 254 414 412 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=48150 $D=0
M1260 413 67 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=43520 $D=0
M1261 414 67 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=48150 $D=0
M1262 9 68 415 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=43520 $D=0
M1263 9 68 416 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=48150 $D=0
M1264 417 69 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=43520 $D=0
M1265 418 69 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=48150 $D=0
M1266 419 415 239 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=43520 $D=0
M1267 420 416 240 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=48150 $D=0
M1268 9 419 749 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=43520 $D=0
M1269 9 420 750 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=48150 $D=0
M1270 421 749 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=43520 $D=0
M1271 422 750 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=48150 $D=0
M1272 419 68 421 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=43520 $D=0
M1273 420 68 422 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=48150 $D=0
M1274 421 417 249 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=43520 $D=0
M1275 422 418 250 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=48150 $D=0
M1276 253 423 421 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=43520 $D=0
M1277 254 424 422 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=48150 $D=0
M1278 423 70 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=43520 $D=0
M1279 424 70 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=48150 $D=0
M1280 9 71 425 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=43520 $D=0
M1281 9 71 426 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=48150 $D=0
M1282 427 72 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=43520 $D=0
M1283 428 72 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=48150 $D=0
M1284 429 425 239 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=43520 $D=0
M1285 430 426 240 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=48150 $D=0
M1286 9 429 751 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=43520 $D=0
M1287 9 430 752 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=48150 $D=0
M1288 431 751 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=43520 $D=0
M1289 432 752 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=48150 $D=0
M1290 429 71 431 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=43520 $D=0
M1291 430 71 432 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=48150 $D=0
M1292 431 427 249 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=43520 $D=0
M1293 432 428 250 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=48150 $D=0
M1294 253 433 431 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=43520 $D=0
M1295 254 434 432 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=48150 $D=0
M1296 433 73 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=43520 $D=0
M1297 434 73 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=48150 $D=0
M1298 9 74 435 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=43520 $D=0
M1299 9 74 436 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=48150 $D=0
M1300 437 75 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=43520 $D=0
M1301 438 75 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=48150 $D=0
M1302 439 435 239 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=43520 $D=0
M1303 440 436 240 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=48150 $D=0
M1304 9 439 753 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=43520 $D=0
M1305 9 440 754 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=48150 $D=0
M1306 441 753 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=43520 $D=0
M1307 442 754 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=48150 $D=0
M1308 439 74 441 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=43520 $D=0
M1309 440 74 442 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=48150 $D=0
M1310 441 437 249 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=43520 $D=0
M1311 442 438 250 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=48150 $D=0
M1312 253 443 441 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=43520 $D=0
M1313 254 444 442 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=48150 $D=0
M1314 443 76 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=43520 $D=0
M1315 444 76 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=48150 $D=0
M1316 9 77 445 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=43520 $D=0
M1317 9 77 446 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=48150 $D=0
M1318 447 78 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=43520 $D=0
M1319 448 78 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=48150 $D=0
M1320 449 445 239 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=43520 $D=0
M1321 450 446 240 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=48150 $D=0
M1322 9 449 755 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=43520 $D=0
M1323 9 450 756 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=48150 $D=0
M1324 451 755 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=43520 $D=0
M1325 452 756 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=48150 $D=0
M1326 449 77 451 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=43520 $D=0
M1327 450 77 452 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=48150 $D=0
M1328 451 447 249 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=43520 $D=0
M1329 452 448 250 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=48150 $D=0
M1330 253 453 451 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=43520 $D=0
M1331 254 454 452 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=48150 $D=0
M1332 453 79 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=43520 $D=0
M1333 454 79 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=48150 $D=0
M1334 9 80 455 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=43520 $D=0
M1335 9 80 456 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=48150 $D=0
M1336 457 81 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=43520 $D=0
M1337 458 81 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=48150 $D=0
M1338 459 455 239 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=43520 $D=0
M1339 460 456 240 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=48150 $D=0
M1340 9 459 757 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=43520 $D=0
M1341 9 460 758 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=48150 $D=0
M1342 461 757 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=43520 $D=0
M1343 462 758 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=48150 $D=0
M1344 459 80 461 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=43520 $D=0
M1345 460 80 462 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=48150 $D=0
M1346 461 457 249 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=43520 $D=0
M1347 462 458 250 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=48150 $D=0
M1348 253 463 461 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=43520 $D=0
M1349 254 464 462 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=48150 $D=0
M1350 463 82 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=43520 $D=0
M1351 464 82 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=48150 $D=0
M1352 9 83 465 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=43520 $D=0
M1353 9 83 466 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=48150 $D=0
M1354 467 84 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=43520 $D=0
M1355 468 84 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=48150 $D=0
M1356 469 465 239 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=43520 $D=0
M1357 470 466 240 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=48150 $D=0
M1358 9 469 759 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=43520 $D=0
M1359 9 470 760 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=48150 $D=0
M1360 471 759 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=43520 $D=0
M1361 472 760 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=48150 $D=0
M1362 469 83 471 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=43520 $D=0
M1363 470 83 472 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=48150 $D=0
M1364 471 467 249 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=43520 $D=0
M1365 472 468 250 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=48150 $D=0
M1366 253 473 471 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=43520 $D=0
M1367 254 474 472 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=48150 $D=0
M1368 473 85 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=43520 $D=0
M1369 474 85 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=48150 $D=0
M1370 9 86 475 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=43520 $D=0
M1371 9 86 476 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=48150 $D=0
M1372 477 87 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=43520 $D=0
M1373 478 87 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=48150 $D=0
M1374 479 475 239 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=43520 $D=0
M1375 480 476 240 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=48150 $D=0
M1376 9 479 761 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=43520 $D=0
M1377 9 480 762 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=48150 $D=0
M1378 481 761 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=43520 $D=0
M1379 482 762 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=48150 $D=0
M1380 479 86 481 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=43520 $D=0
M1381 480 86 482 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=48150 $D=0
M1382 481 477 249 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=43520 $D=0
M1383 482 478 250 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=48150 $D=0
M1384 253 483 481 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=43520 $D=0
M1385 254 484 482 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=48150 $D=0
M1386 483 88 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=43520 $D=0
M1387 484 88 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=48150 $D=0
M1388 9 89 485 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=43520 $D=0
M1389 9 89 486 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=48150 $D=0
M1390 487 90 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=43520 $D=0
M1391 488 90 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=48150 $D=0
M1392 489 485 239 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=43520 $D=0
M1393 490 486 240 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=48150 $D=0
M1394 9 489 763 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=43520 $D=0
M1395 9 490 764 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=48150 $D=0
M1396 491 763 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=43520 $D=0
M1397 492 764 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=48150 $D=0
M1398 489 89 491 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=43520 $D=0
M1399 490 89 492 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=48150 $D=0
M1400 491 487 249 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=43520 $D=0
M1401 492 488 250 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=48150 $D=0
M1402 253 493 491 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=43520 $D=0
M1403 254 494 492 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=48150 $D=0
M1404 493 91 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=43520 $D=0
M1405 494 91 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=48150 $D=0
M1406 9 92 495 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=43520 $D=0
M1407 9 92 496 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=48150 $D=0
M1408 497 93 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=43520 $D=0
M1409 498 93 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=48150 $D=0
M1410 499 495 239 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=43520 $D=0
M1411 500 496 240 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=48150 $D=0
M1412 9 499 765 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=43520 $D=0
M1413 9 500 766 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=48150 $D=0
M1414 501 765 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=43520 $D=0
M1415 502 766 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=48150 $D=0
M1416 499 92 501 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=43520 $D=0
M1417 500 92 502 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=48150 $D=0
M1418 501 497 249 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=43520 $D=0
M1419 502 498 250 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=48150 $D=0
M1420 253 503 501 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=43520 $D=0
M1421 254 504 502 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=48150 $D=0
M1422 503 94 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=43520 $D=0
M1423 504 94 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=48150 $D=0
M1424 9 95 505 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=43520 $D=0
M1425 9 95 506 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=48150 $D=0
M1426 507 96 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=43520 $D=0
M1427 508 96 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=48150 $D=0
M1428 509 505 239 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=43520 $D=0
M1429 510 506 240 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=48150 $D=0
M1430 9 509 767 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=43520 $D=0
M1431 9 510 768 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=48150 $D=0
M1432 511 767 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=43520 $D=0
M1433 512 768 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=48150 $D=0
M1434 509 95 511 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=43520 $D=0
M1435 510 95 512 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=48150 $D=0
M1436 511 507 249 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=43520 $D=0
M1437 512 508 250 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=48150 $D=0
M1438 253 513 511 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=43520 $D=0
M1439 254 514 512 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=48150 $D=0
M1440 513 97 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=43520 $D=0
M1441 514 97 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=48150 $D=0
M1442 9 98 515 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=43520 $D=0
M1443 9 98 516 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=48150 $D=0
M1444 517 99 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=43520 $D=0
M1445 518 99 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=48150 $D=0
M1446 519 515 239 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=43520 $D=0
M1447 520 516 240 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=48150 $D=0
M1448 9 519 769 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=43520 $D=0
M1449 9 520 770 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=48150 $D=0
M1450 521 769 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=43520 $D=0
M1451 522 770 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=48150 $D=0
M1452 519 98 521 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=43520 $D=0
M1453 520 98 522 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=48150 $D=0
M1454 521 517 249 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=43520 $D=0
M1455 522 518 250 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=48150 $D=0
M1456 253 523 521 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=43520 $D=0
M1457 254 524 522 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=48150 $D=0
M1458 523 100 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=43520 $D=0
M1459 524 100 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=48150 $D=0
M1460 9 101 525 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=43520 $D=0
M1461 9 101 526 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=48150 $D=0
M1462 527 102 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=43520 $D=0
M1463 528 102 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=48150 $D=0
M1464 529 525 239 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=43520 $D=0
M1465 530 526 240 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=48150 $D=0
M1466 9 529 771 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=43520 $D=0
M1467 9 530 772 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=48150 $D=0
M1468 531 771 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=43520 $D=0
M1469 532 772 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=48150 $D=0
M1470 529 101 531 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=43520 $D=0
M1471 530 101 532 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=48150 $D=0
M1472 531 527 249 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=43520 $D=0
M1473 532 528 250 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=48150 $D=0
M1474 253 533 531 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=43520 $D=0
M1475 254 534 532 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=48150 $D=0
M1476 533 103 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=43520 $D=0
M1477 534 103 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=48150 $D=0
M1478 9 104 535 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=43520 $D=0
M1479 9 104 536 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=48150 $D=0
M1480 537 105 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=43520 $D=0
M1481 538 105 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=48150 $D=0
M1482 539 535 239 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=43520 $D=0
M1483 540 536 240 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=48150 $D=0
M1484 9 539 773 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=43520 $D=0
M1485 9 540 774 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=48150 $D=0
M1486 541 773 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=43520 $D=0
M1487 542 774 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=48150 $D=0
M1488 539 104 541 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=43520 $D=0
M1489 540 104 542 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=48150 $D=0
M1490 541 537 249 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=43520 $D=0
M1491 542 538 250 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=48150 $D=0
M1492 253 543 541 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=43520 $D=0
M1493 254 544 542 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=48150 $D=0
M1494 543 109 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=43520 $D=0
M1495 544 109 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=48150 $D=0
M1496 9 110 545 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=43520 $D=0
M1497 9 110 546 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=48150 $D=0
M1498 547 111 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=43520 $D=0
M1499 548 111 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=48150 $D=0
M1500 549 545 239 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=43520 $D=0
M1501 550 546 240 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=48150 $D=0
M1502 9 549 775 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=43520 $D=0
M1503 9 550 776 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=48150 $D=0
M1504 551 775 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=43520 $D=0
M1505 552 776 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=48150 $D=0
M1506 549 110 551 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=43520 $D=0
M1507 550 110 552 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=48150 $D=0
M1508 551 547 249 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=43520 $D=0
M1509 552 548 250 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=48150 $D=0
M1510 253 553 551 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=43520 $D=0
M1511 254 554 552 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=48150 $D=0
M1512 553 113 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=43520 $D=0
M1513 554 113 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=48150 $D=0
M1514 9 114 555 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=43520 $D=0
M1515 9 114 556 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=48150 $D=0
M1516 557 115 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=43520 $D=0
M1517 558 115 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=48150 $D=0
M1518 6 557 249 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=43520 $D=0
M1519 6 558 250 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=48150 $D=0
M1520 253 555 6 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=43520 $D=0
M1521 254 556 6 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=48150 $D=0
M1522 9 561 559 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=43520 $D=0
M1523 9 562 560 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=48150 $D=0
M1524 561 117 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=43520 $D=0
M1525 562 117 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=48150 $D=0
M1526 777 249 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=43520 $D=0
M1527 778 250 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=48150 $D=0
M1528 563 561 777 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=43520 $D=0
M1529 564 562 778 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=48150 $D=0
M1530 9 563 565 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=43520 $D=0
M1531 9 564 566 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=48150 $D=0
M1532 779 565 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=43520 $D=0
M1533 780 566 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=48150 $D=0
M1534 563 559 779 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=43520 $D=0
M1535 564 560 780 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=48150 $D=0
M1536 9 569 567 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=43520 $D=0
M1537 9 570 568 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=48150 $D=0
M1538 569 117 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=43520 $D=0
M1539 570 117 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=48150 $D=0
M1540 781 253 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=43520 $D=0
M1541 782 254 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=48150 $D=0
M1542 571 569 781 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=43520 $D=0
M1543 572 570 782 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=48150 $D=0
M1544 9 571 119 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=43520 $D=0
M1545 9 572 120 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=48150 $D=0
M1546 783 119 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=43520 $D=0
M1547 784 120 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=48150 $D=0
M1548 571 567 783 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=43520 $D=0
M1549 572 568 784 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=48150 $D=0
M1550 573 121 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=43520 $D=0
M1551 574 121 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=48150 $D=0
M1552 575 121 565 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=43520 $D=0
M1553 576 121 566 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=48150 $D=0
M1554 122 573 575 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=43520 $D=0
M1555 123 574 576 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=48150 $D=0
M1556 577 124 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=43520 $D=0
M1557 578 124 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=48150 $D=0
M1558 579 124 119 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=43520 $D=0
M1559 580 124 120 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=48150 $D=0
M1560 785 577 579 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=43520 $D=0
M1561 786 578 580 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=48150 $D=0
M1562 9 119 785 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=43520 $D=0
M1563 9 120 786 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=48150 $D=0
M1564 581 125 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=43520 $D=0
M1565 582 125 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=48150 $D=0
M1566 583 125 579 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=43520 $D=0
M1567 584 125 580 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=48150 $D=0
M1568 11 581 583 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=43520 $D=0
M1569 12 582 584 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=48150 $D=0
M1570 586 585 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=43520 $D=0
M1571 587 126 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=48150 $D=0
M1572 9 590 588 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=43520 $D=0
M1573 9 591 589 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=48150 $D=0
M1574 592 575 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=43520 $D=0
M1575 593 576 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=48150 $D=0
M1576 590 575 585 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=43520 $D=0
M1577 591 576 126 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=48150 $D=0
M1578 586 592 590 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=43520 $D=0
M1579 587 593 591 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=48150 $D=0
M1580 594 588 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=43520 $D=0
M1581 595 589 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=48150 $D=0
M1582 127 588 583 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=43520 $D=0
M1583 585 589 584 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=48150 $D=0
M1584 575 594 127 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=43520 $D=0
M1585 576 595 585 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=48150 $D=0
M1586 596 127 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=43520 $D=0
M1587 597 585 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=48150 $D=0
M1588 598 588 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=43520 $D=0
M1589 599 589 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=48150 $D=0
M1590 600 588 596 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=43520 $D=0
M1591 601 589 597 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=48150 $D=0
M1592 583 598 600 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=43520 $D=0
M1593 584 599 601 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=48150 $D=0
M1594 797 575 9 9 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=43160 $D=0
M1595 798 576 9 9 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=47790 $D=0
M1596 602 583 797 9 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=43160 $D=0
M1597 603 584 798 9 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=47790 $D=0
M1598 604 600 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=43520 $D=0
M1599 605 601 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=48150 $D=0
M1600 606 575 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=43520 $D=0
M1601 607 576 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=48150 $D=0
M1602 9 583 606 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=43520 $D=0
M1603 9 584 607 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=48150 $D=0
M1604 608 575 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=43520 $D=0
M1605 609 576 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=48150 $D=0
M1606 9 583 608 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=43520 $D=0
M1607 9 584 609 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=48150 $D=0
M1608 799 575 9 9 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=43340 $D=0
M1609 800 576 9 9 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=47970 $D=0
M1610 612 583 799 9 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=43340 $D=0
M1611 613 584 800 9 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=47970 $D=0
M1612 9 608 612 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=43520 $D=0
M1613 9 609 613 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=48150 $D=0
M1614 614 130 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=43520 $D=0
M1615 615 130 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=48150 $D=0
M1616 616 130 602 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=43520 $D=0
M1617 617 130 603 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=48150 $D=0
M1618 606 614 616 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=43520 $D=0
M1619 607 615 617 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=48150 $D=0
M1620 618 130 604 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=43520 $D=0
M1621 619 130 605 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=48150 $D=0
M1622 612 614 618 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=43520 $D=0
M1623 613 615 619 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=48150 $D=0
M1624 620 131 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=43520 $D=0
M1625 621 131 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=48150 $D=0
M1626 622 131 618 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=43520 $D=0
M1627 623 131 619 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=48150 $D=0
M1628 616 620 622 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=43520 $D=0
M1629 617 621 623 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=48150 $D=0
M1630 13 622 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=43520 $D=0
M1631 14 623 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=48150 $D=0
M1632 624 132 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=43520 $D=0
M1633 625 132 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=48150 $D=0
M1634 626 132 133 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=43520 $D=0
M1635 627 132 134 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=48150 $D=0
M1636 135 624 626 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=43520 $D=0
M1637 136 625 627 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=48150 $D=0
M1638 628 132 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=43520 $D=0
M1639 629 132 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=48150 $D=0
M1640 630 132 137 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=43520 $D=0
M1641 631 132 138 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=48150 $D=0
M1642 139 628 630 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=43520 $D=0
M1643 140 629 631 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=48150 $D=0
M1644 632 132 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=43520 $D=0
M1645 633 132 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=48150 $D=0
M1646 634 132 129 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=43520 $D=0
M1647 635 132 128 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=48150 $D=0
M1648 141 632 634 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=43520 $D=0
M1649 108 633 635 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=48150 $D=0
M1650 636 132 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=43520 $D=0
M1651 637 132 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=48150 $D=0
M1652 638 132 142 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=43520 $D=0
M1653 639 132 143 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=48150 $D=0
M1654 144 636 638 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=43520 $D=0
M1655 145 637 639 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=48150 $D=0
M1656 640 132 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=43520 $D=0
M1657 641 132 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=48150 $D=0
M1658 642 132 146 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=43520 $D=0
M1659 643 132 147 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=48150 $D=0
M1660 148 640 642 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=43520 $D=0
M1661 148 641 643 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=48150 $D=0
M1662 9 575 787 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=43520 $D=0
M1663 9 576 788 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=48150 $D=0
M1664 136 787 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=43520 $D=0
M1665 133 788 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=48150 $D=0
M1666 644 149 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=43520 $D=0
M1667 645 149 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=48150 $D=0
M1668 150 149 136 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=43520 $D=0
M1669 151 149 133 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=48150 $D=0
M1670 626 644 150 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=43520 $D=0
M1671 627 645 151 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=48150 $D=0
M1672 646 152 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=43520 $D=0
M1673 647 152 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=48150 $D=0
M1674 153 152 150 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=43520 $D=0
M1675 116 152 151 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=48150 $D=0
M1676 630 646 153 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=43520 $D=0
M1677 631 647 116 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=48150 $D=0
M1678 648 154 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=43520 $D=0
M1679 649 154 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=48150 $D=0
M1680 155 154 153 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=43520 $D=0
M1681 106 154 116 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=48150 $D=0
M1682 634 648 155 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=43520 $D=0
M1683 635 649 106 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=48150 $D=0
M1684 650 156 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=43520 $D=0
M1685 651 156 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=48150 $D=0
M1686 157 156 155 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=43520 $D=0
M1687 158 156 106 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=48150 $D=0
M1688 638 650 157 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=43520 $D=0
M1689 639 651 158 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=48150 $D=0
M1690 652 159 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=43520 $D=0
M1691 653 159 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=48150 $D=0
M1692 225 159 157 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=43520 $D=0
M1693 226 159 158 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=48150 $D=0
M1694 642 652 225 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=43520 $D=0
M1695 643 653 226 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=48150 $D=0
M1696 654 160 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=43520 $D=0
M1697 655 160 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=48150 $D=0
M1698 656 160 119 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=43520 $D=0
M1699 657 160 120 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=48150 $D=0
M1700 11 654 656 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=43520 $D=0
M1701 12 655 657 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=48150 $D=0
M1702 658 565 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=43520 $D=0
M1703 659 566 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=48150 $D=0
M1704 9 656 658 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=43520 $D=0
M1705 9 657 659 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=48150 $D=0
M1706 801 565 9 9 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=43340 $D=0
M1707 802 566 9 9 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=47970 $D=0
M1708 662 656 801 9 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=43340 $D=0
M1709 663 657 802 9 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=47970 $D=0
M1710 9 658 662 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=43520 $D=0
M1711 9 659 663 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=48150 $D=0
M1712 789 161 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=43520 $D=0
M1713 790 664 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=48150 $D=0
M1714 9 662 789 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=43520 $D=0
M1715 9 663 790 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=48150 $D=0
M1716 664 789 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=43520 $D=0
M1717 162 790 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=48150 $D=0
M1718 803 565 9 9 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=43160 $D=0
M1719 804 566 9 9 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=47790 $D=0
M1720 665 667 803 9 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=43160 $D=0
M1721 666 668 804 9 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=47790 $D=0
M1722 667 656 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=43520 $D=0
M1723 668 657 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=48150 $D=0
M1724 669 665 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=43520 $D=0
M1725 670 666 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=48150 $D=0
M1726 9 161 669 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=43520 $D=0
M1727 9 664 670 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=48150 $D=0
M1728 672 163 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=43520 $D=0
M1729 673 671 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=48150 $D=0
M1730 671 669 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=43520 $D=0
M1731 164 670 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=48150 $D=0
M1732 9 672 671 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=43520 $D=0
M1733 9 673 164 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=48150 $D=0
M1734 675 674 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=43520 $D=0
M1735 676 165 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=48150 $D=0
M1736 9 679 677 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=43520 $D=0
M1737 9 680 678 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=48150 $D=0
M1738 681 122 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=43520 $D=0
M1739 682 123 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=48150 $D=0
M1740 679 122 674 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=43520 $D=0
M1741 680 123 165 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=48150 $D=0
M1742 675 681 679 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=43520 $D=0
M1743 676 682 680 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=48150 $D=0
M1744 683 677 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=43520 $D=0
M1745 684 678 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=48150 $D=0
M1746 166 677 6 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=43520 $D=0
M1747 674 678 6 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=48150 $D=0
M1748 122 683 166 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=43520 $D=0
M1749 123 684 674 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=48150 $D=0
M1750 685 166 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=43520 $D=0
M1751 686 674 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=48150 $D=0
M1752 687 677 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=43520 $D=0
M1753 688 678 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=48150 $D=0
M1754 227 677 685 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=43520 $D=0
M1755 228 678 686 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=48150 $D=0
M1756 6 687 227 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=43520 $D=0
M1757 6 688 228 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=48150 $D=0
M1758 689 167 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=43520 $D=0
M1759 690 167 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=48150 $D=0
M1760 691 167 227 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=43520 $D=0
M1761 692 167 228 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=48150 $D=0
M1762 13 689 691 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=43520 $D=0
M1763 14 690 692 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=48150 $D=0
M1764 693 168 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=43520 $D=0
M1765 694 168 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=48150 $D=0
M1766 695 168 691 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=43520 $D=0
M1767 696 168 692 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=48150 $D=0
M1768 6 693 695 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=43520 $D=0
M1769 6 694 696 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=48150 $D=0
M1770 697 117 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=43520 $D=0
M1771 698 117 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=48150 $D=0
M1772 9 697 699 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=43520 $D=0
M1773 9 698 700 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=48150 $D=0
M1774 701 117 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=43520 $D=0
M1775 702 117 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=48150 $D=0
M1776 703 699 695 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=43520 $D=0
M1777 704 700 696 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=48150 $D=0
M1778 9 703 791 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=43520 $D=0
M1779 9 704 792 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=48150 $D=0
M1780 705 791 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=43520 $D=0
M1781 706 792 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=48150 $D=0
M1782 703 697 705 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=43520 $D=0
M1783 704 698 706 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=48150 $D=0
M1784 707 701 705 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=43520 $D=0
M1785 708 702 706 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=48150 $D=0
M1786 9 711 709 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=43520 $D=0
M1787 9 712 710 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=48150 $D=0
M1788 711 117 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=43520 $D=0
M1789 712 117 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=48150 $D=0
M1790 793 707 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=43520 $D=0
M1791 794 708 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=48150 $D=0
M1792 713 711 793 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=43520 $D=0
M1793 714 712 794 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=48150 $D=0
M1794 9 713 122 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=43520 $D=0
M1795 9 714 123 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=48150 $D=0
M1796 795 122 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=43520 $D=0
M1797 796 123 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=48150 $D=0
M1798 713 709 795 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=43520 $D=0
M1799 714 710 796 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=48150 $D=0
.ENDS
***************************************
.SUBCKT ICV_38 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 108 109 111 112 113 115 116 117 118 119 120 121 122 123
+ 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141 142 143
+ 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162 163
+ 164 165 166 167
** N=811 EP=164 IP=1514 FDC=1800
M0 196 1 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=33010 $D=1
M1 197 1 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=37640 $D=1
M2 198 196 2 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=33010 $D=1
M3 199 197 3 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=37640 $D=1
M4 6 1 198 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=33010 $D=1
M5 6 1 199 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=37640 $D=1
M6 200 196 4 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=33010 $D=1
M7 201 197 4 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=37640 $D=1
M8 5 1 200 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=33010 $D=1
M9 5 1 201 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=37640 $D=1
M10 202 196 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=33010 $D=1
M11 203 197 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=37640 $D=1
M12 6 1 202 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=33010 $D=1
M13 6 1 203 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=37640 $D=1
M14 206 204 202 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=33010 $D=1
M15 207 205 203 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=37640 $D=1
M16 204 7 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=33010 $D=1
M17 205 7 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=37640 $D=1
M18 208 204 200 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=33010 $D=1
M19 209 205 201 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=37640 $D=1
M20 198 7 208 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=33010 $D=1
M21 199 7 209 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=37640 $D=1
M22 210 8 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=33010 $D=1
M23 211 8 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=37640 $D=1
M24 212 210 208 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=33010 $D=1
M25 213 211 209 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=37640 $D=1
M26 206 8 212 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=33010 $D=1
M27 207 8 213 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=37640 $D=1
M28 214 10 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=33010 $D=1
M29 215 10 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=37640 $D=1
M30 216 214 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=33010 $D=1
M31 217 215 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=37640 $D=1
M32 11 10 216 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=33010 $D=1
M33 12 10 217 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=37640 $D=1
M34 218 214 13 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=33010 $D=1
M35 219 215 14 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=37640 $D=1
M36 220 10 218 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=33010 $D=1
M37 221 10 219 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=37640 $D=1
M38 224 214 222 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=33010 $D=1
M39 225 215 223 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=37640 $D=1
M40 212 10 224 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=33010 $D=1
M41 213 10 225 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=37640 $D=1
M42 228 226 224 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=33010 $D=1
M43 229 227 225 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=37640 $D=1
M44 226 15 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=33010 $D=1
M45 227 15 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=37640 $D=1
M46 230 226 218 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=33010 $D=1
M47 231 227 219 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=37640 $D=1
M48 216 15 230 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=33010 $D=1
M49 217 15 231 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=37640 $D=1
M50 232 16 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=33010 $D=1
M51 233 16 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=37640 $D=1
M52 234 232 230 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=33010 $D=1
M53 235 233 231 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=37640 $D=1
M54 228 16 234 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=33010 $D=1
M55 229 16 235 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=37640 $D=1
M56 6 17 236 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=33010 $D=1
M57 6 17 237 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=37640 $D=1
M58 238 18 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=33010 $D=1
M59 239 18 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=37640 $D=1
M60 240 17 234 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=33010 $D=1
M61 241 17 235 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=37640 $D=1
M62 6 240 710 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=33010 $D=1
M63 6 241 711 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=37640 $D=1
M64 242 710 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=33010 $D=1
M65 243 711 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=37640 $D=1
M66 240 236 242 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=33010 $D=1
M67 241 237 243 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=37640 $D=1
M68 242 18 244 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=33010 $D=1
M69 243 18 245 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=37640 $D=1
M70 248 19 242 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=33010 $D=1
M71 249 19 243 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=37640 $D=1
M72 246 19 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=33010 $D=1
M73 247 19 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=37640 $D=1
M74 6 20 250 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=33010 $D=1
M75 6 20 251 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=37640 $D=1
M76 252 21 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=33010 $D=1
M77 253 21 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=37640 $D=1
M78 254 20 234 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=33010 $D=1
M79 255 20 235 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=37640 $D=1
M80 6 254 712 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=33010 $D=1
M81 6 255 713 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=37640 $D=1
M82 256 712 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=33010 $D=1
M83 257 713 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=37640 $D=1
M84 254 250 256 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=33010 $D=1
M85 255 251 257 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=37640 $D=1
M86 256 21 244 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=33010 $D=1
M87 257 21 245 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=37640 $D=1
M88 248 22 256 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=33010 $D=1
M89 249 22 257 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=37640 $D=1
M90 258 22 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=33010 $D=1
M91 259 22 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=37640 $D=1
M92 6 23 260 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=33010 $D=1
M93 6 23 261 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=37640 $D=1
M94 262 24 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=33010 $D=1
M95 263 24 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=37640 $D=1
M96 264 23 234 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=33010 $D=1
M97 265 23 235 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=37640 $D=1
M98 6 264 714 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=33010 $D=1
M99 6 265 715 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=37640 $D=1
M100 266 714 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=33010 $D=1
M101 267 715 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=37640 $D=1
M102 264 260 266 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=33010 $D=1
M103 265 261 267 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=37640 $D=1
M104 266 24 244 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=33010 $D=1
M105 267 24 245 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=37640 $D=1
M106 248 25 266 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=33010 $D=1
M107 249 25 267 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=37640 $D=1
M108 268 25 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=33010 $D=1
M109 269 25 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=37640 $D=1
M110 6 26 270 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=33010 $D=1
M111 6 26 271 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=37640 $D=1
M112 272 27 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=33010 $D=1
M113 273 27 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=37640 $D=1
M114 274 26 234 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=33010 $D=1
M115 275 26 235 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=37640 $D=1
M116 6 274 716 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=33010 $D=1
M117 6 275 717 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=37640 $D=1
M118 276 716 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=33010 $D=1
M119 277 717 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=37640 $D=1
M120 274 270 276 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=33010 $D=1
M121 275 271 277 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=37640 $D=1
M122 276 27 244 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=33010 $D=1
M123 277 27 245 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=37640 $D=1
M124 248 28 276 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=33010 $D=1
M125 249 28 277 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=37640 $D=1
M126 278 28 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=33010 $D=1
M127 279 28 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=37640 $D=1
M128 6 29 280 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=33010 $D=1
M129 6 29 281 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=37640 $D=1
M130 282 30 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=33010 $D=1
M131 283 30 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=37640 $D=1
M132 284 29 234 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=33010 $D=1
M133 285 29 235 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=37640 $D=1
M134 6 284 718 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=33010 $D=1
M135 6 285 719 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=37640 $D=1
M136 286 718 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=33010 $D=1
M137 287 719 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=37640 $D=1
M138 284 280 286 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=33010 $D=1
M139 285 281 287 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=37640 $D=1
M140 286 30 244 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=33010 $D=1
M141 287 30 245 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=37640 $D=1
M142 248 31 286 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=33010 $D=1
M143 249 31 287 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=37640 $D=1
M144 288 31 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=33010 $D=1
M145 289 31 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=37640 $D=1
M146 6 32 290 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=33010 $D=1
M147 6 32 291 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=37640 $D=1
M148 292 33 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=33010 $D=1
M149 293 33 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=37640 $D=1
M150 294 32 234 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=33010 $D=1
M151 295 32 235 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=37640 $D=1
M152 6 294 720 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=33010 $D=1
M153 6 295 721 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=37640 $D=1
M154 296 720 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=33010 $D=1
M155 297 721 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=37640 $D=1
M156 294 290 296 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=33010 $D=1
M157 295 291 297 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=37640 $D=1
M158 296 33 244 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=33010 $D=1
M159 297 33 245 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=37640 $D=1
M160 248 34 296 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=33010 $D=1
M161 249 34 297 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=37640 $D=1
M162 298 34 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=33010 $D=1
M163 299 34 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=37640 $D=1
M164 6 35 300 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=33010 $D=1
M165 6 35 301 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=37640 $D=1
M166 302 36 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=33010 $D=1
M167 303 36 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=37640 $D=1
M168 304 35 234 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=33010 $D=1
M169 305 35 235 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=37640 $D=1
M170 6 304 722 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=33010 $D=1
M171 6 305 723 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=37640 $D=1
M172 306 722 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=33010 $D=1
M173 307 723 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=37640 $D=1
M174 304 300 306 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=33010 $D=1
M175 305 301 307 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=37640 $D=1
M176 306 36 244 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=33010 $D=1
M177 307 36 245 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=37640 $D=1
M178 248 37 306 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=33010 $D=1
M179 249 37 307 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=37640 $D=1
M180 308 37 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=33010 $D=1
M181 309 37 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=37640 $D=1
M182 6 38 310 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=33010 $D=1
M183 6 38 311 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=37640 $D=1
M184 312 39 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=33010 $D=1
M185 313 39 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=37640 $D=1
M186 314 38 234 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=33010 $D=1
M187 315 38 235 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=37640 $D=1
M188 6 314 724 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=33010 $D=1
M189 6 315 725 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=37640 $D=1
M190 316 724 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=33010 $D=1
M191 317 725 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=37640 $D=1
M192 314 310 316 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=33010 $D=1
M193 315 311 317 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=37640 $D=1
M194 316 39 244 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=33010 $D=1
M195 317 39 245 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=37640 $D=1
M196 248 40 316 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=33010 $D=1
M197 249 40 317 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=37640 $D=1
M198 318 40 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=33010 $D=1
M199 319 40 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=37640 $D=1
M200 6 41 320 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=33010 $D=1
M201 6 41 321 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=37640 $D=1
M202 322 42 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=33010 $D=1
M203 323 42 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=37640 $D=1
M204 324 41 234 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=33010 $D=1
M205 325 41 235 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=37640 $D=1
M206 6 324 726 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=33010 $D=1
M207 6 325 727 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=37640 $D=1
M208 326 726 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=33010 $D=1
M209 327 727 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=37640 $D=1
M210 324 320 326 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=33010 $D=1
M211 325 321 327 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=37640 $D=1
M212 326 42 244 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=33010 $D=1
M213 327 42 245 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=37640 $D=1
M214 248 43 326 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=33010 $D=1
M215 249 43 327 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=37640 $D=1
M216 328 43 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=33010 $D=1
M217 329 43 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=37640 $D=1
M218 6 44 330 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=33010 $D=1
M219 6 44 331 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=37640 $D=1
M220 332 45 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=33010 $D=1
M221 333 45 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=37640 $D=1
M222 334 44 234 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=33010 $D=1
M223 335 44 235 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=37640 $D=1
M224 6 334 728 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=33010 $D=1
M225 6 335 729 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=37640 $D=1
M226 336 728 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=33010 $D=1
M227 337 729 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=37640 $D=1
M228 334 330 336 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=33010 $D=1
M229 335 331 337 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=37640 $D=1
M230 336 45 244 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=33010 $D=1
M231 337 45 245 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=37640 $D=1
M232 248 46 336 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=33010 $D=1
M233 249 46 337 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=37640 $D=1
M234 338 46 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=33010 $D=1
M235 339 46 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=37640 $D=1
M236 6 47 340 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=33010 $D=1
M237 6 47 341 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=37640 $D=1
M238 342 48 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=33010 $D=1
M239 343 48 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=37640 $D=1
M240 344 47 234 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=33010 $D=1
M241 345 47 235 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=37640 $D=1
M242 6 344 730 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=33010 $D=1
M243 6 345 731 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=37640 $D=1
M244 346 730 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=33010 $D=1
M245 347 731 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=37640 $D=1
M246 344 340 346 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=33010 $D=1
M247 345 341 347 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=37640 $D=1
M248 346 48 244 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=33010 $D=1
M249 347 48 245 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=37640 $D=1
M250 248 49 346 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=33010 $D=1
M251 249 49 347 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=37640 $D=1
M252 348 49 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=33010 $D=1
M253 349 49 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=37640 $D=1
M254 6 50 350 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=33010 $D=1
M255 6 50 351 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=37640 $D=1
M256 352 51 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=33010 $D=1
M257 353 51 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=37640 $D=1
M258 354 50 234 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=33010 $D=1
M259 355 50 235 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=37640 $D=1
M260 6 354 732 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=33010 $D=1
M261 6 355 733 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=37640 $D=1
M262 356 732 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=33010 $D=1
M263 357 733 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=37640 $D=1
M264 354 350 356 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=33010 $D=1
M265 355 351 357 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=37640 $D=1
M266 356 51 244 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=33010 $D=1
M267 357 51 245 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=37640 $D=1
M268 248 52 356 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=33010 $D=1
M269 249 52 357 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=37640 $D=1
M270 358 52 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=33010 $D=1
M271 359 52 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=37640 $D=1
M272 6 53 360 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=33010 $D=1
M273 6 53 361 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=37640 $D=1
M274 362 54 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=33010 $D=1
M275 363 54 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=37640 $D=1
M276 364 53 234 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=33010 $D=1
M277 365 53 235 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=37640 $D=1
M278 6 364 734 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=33010 $D=1
M279 6 365 735 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=37640 $D=1
M280 366 734 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=33010 $D=1
M281 367 735 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=37640 $D=1
M282 364 360 366 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=33010 $D=1
M283 365 361 367 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=37640 $D=1
M284 366 54 244 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=33010 $D=1
M285 367 54 245 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=37640 $D=1
M286 248 55 366 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=33010 $D=1
M287 249 55 367 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=37640 $D=1
M288 368 55 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=33010 $D=1
M289 369 55 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=37640 $D=1
M290 6 56 370 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=33010 $D=1
M291 6 56 371 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=37640 $D=1
M292 372 57 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=33010 $D=1
M293 373 57 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=37640 $D=1
M294 374 56 234 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=33010 $D=1
M295 375 56 235 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=37640 $D=1
M296 6 374 736 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=33010 $D=1
M297 6 375 737 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=37640 $D=1
M298 376 736 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=33010 $D=1
M299 377 737 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=37640 $D=1
M300 374 370 376 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=33010 $D=1
M301 375 371 377 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=37640 $D=1
M302 376 57 244 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=33010 $D=1
M303 377 57 245 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=37640 $D=1
M304 248 58 376 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=33010 $D=1
M305 249 58 377 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=37640 $D=1
M306 378 58 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=33010 $D=1
M307 379 58 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=37640 $D=1
M308 6 59 380 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=33010 $D=1
M309 6 59 381 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=37640 $D=1
M310 382 60 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=33010 $D=1
M311 383 60 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=37640 $D=1
M312 384 59 234 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=33010 $D=1
M313 385 59 235 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=37640 $D=1
M314 6 384 738 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=33010 $D=1
M315 6 385 739 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=37640 $D=1
M316 386 738 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=33010 $D=1
M317 387 739 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=37640 $D=1
M318 384 380 386 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=33010 $D=1
M319 385 381 387 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=37640 $D=1
M320 386 60 244 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=33010 $D=1
M321 387 60 245 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=37640 $D=1
M322 248 61 386 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=33010 $D=1
M323 249 61 387 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=37640 $D=1
M324 388 61 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=33010 $D=1
M325 389 61 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=37640 $D=1
M326 6 62 390 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=33010 $D=1
M327 6 62 391 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=37640 $D=1
M328 392 63 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=33010 $D=1
M329 393 63 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=37640 $D=1
M330 394 62 234 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=33010 $D=1
M331 395 62 235 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=37640 $D=1
M332 6 394 740 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=33010 $D=1
M333 6 395 741 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=37640 $D=1
M334 396 740 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=33010 $D=1
M335 397 741 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=37640 $D=1
M336 394 390 396 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=33010 $D=1
M337 395 391 397 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=37640 $D=1
M338 396 63 244 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=33010 $D=1
M339 397 63 245 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=37640 $D=1
M340 248 64 396 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=33010 $D=1
M341 249 64 397 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=37640 $D=1
M342 398 64 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=33010 $D=1
M343 399 64 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=37640 $D=1
M344 6 65 400 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=33010 $D=1
M345 6 65 401 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=37640 $D=1
M346 402 66 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=33010 $D=1
M347 403 66 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=37640 $D=1
M348 404 65 234 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=33010 $D=1
M349 405 65 235 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=37640 $D=1
M350 6 404 742 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=33010 $D=1
M351 6 405 743 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=37640 $D=1
M352 406 742 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=33010 $D=1
M353 407 743 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=37640 $D=1
M354 404 400 406 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=33010 $D=1
M355 405 401 407 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=37640 $D=1
M356 406 66 244 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=33010 $D=1
M357 407 66 245 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=37640 $D=1
M358 248 67 406 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=33010 $D=1
M359 249 67 407 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=37640 $D=1
M360 408 67 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=33010 $D=1
M361 409 67 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=37640 $D=1
M362 6 68 410 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=33010 $D=1
M363 6 68 411 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=37640 $D=1
M364 412 69 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=33010 $D=1
M365 413 69 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=37640 $D=1
M366 414 68 234 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=33010 $D=1
M367 415 68 235 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=37640 $D=1
M368 6 414 744 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=33010 $D=1
M369 6 415 745 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=37640 $D=1
M370 416 744 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=33010 $D=1
M371 417 745 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=37640 $D=1
M372 414 410 416 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=33010 $D=1
M373 415 411 417 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=37640 $D=1
M374 416 69 244 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=33010 $D=1
M375 417 69 245 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=37640 $D=1
M376 248 70 416 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=33010 $D=1
M377 249 70 417 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=37640 $D=1
M378 418 70 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=33010 $D=1
M379 419 70 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=37640 $D=1
M380 6 71 420 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=33010 $D=1
M381 6 71 421 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=37640 $D=1
M382 422 72 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=33010 $D=1
M383 423 72 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=37640 $D=1
M384 424 71 234 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=33010 $D=1
M385 425 71 235 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=37640 $D=1
M386 6 424 746 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=33010 $D=1
M387 6 425 747 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=37640 $D=1
M388 426 746 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=33010 $D=1
M389 427 747 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=37640 $D=1
M390 424 420 426 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=33010 $D=1
M391 425 421 427 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=37640 $D=1
M392 426 72 244 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=33010 $D=1
M393 427 72 245 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=37640 $D=1
M394 248 73 426 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=33010 $D=1
M395 249 73 427 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=37640 $D=1
M396 428 73 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=33010 $D=1
M397 429 73 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=37640 $D=1
M398 6 74 430 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=33010 $D=1
M399 6 74 431 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=37640 $D=1
M400 432 75 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=33010 $D=1
M401 433 75 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=37640 $D=1
M402 434 74 234 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=33010 $D=1
M403 435 74 235 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=37640 $D=1
M404 6 434 748 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=33010 $D=1
M405 6 435 749 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=37640 $D=1
M406 436 748 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=33010 $D=1
M407 437 749 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=37640 $D=1
M408 434 430 436 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=33010 $D=1
M409 435 431 437 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=37640 $D=1
M410 436 75 244 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=33010 $D=1
M411 437 75 245 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=37640 $D=1
M412 248 76 436 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=33010 $D=1
M413 249 76 437 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=37640 $D=1
M414 438 76 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=33010 $D=1
M415 439 76 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=37640 $D=1
M416 6 77 440 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=33010 $D=1
M417 6 77 441 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=37640 $D=1
M418 442 78 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=33010 $D=1
M419 443 78 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=37640 $D=1
M420 444 77 234 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=33010 $D=1
M421 445 77 235 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=37640 $D=1
M422 6 444 750 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=33010 $D=1
M423 6 445 751 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=37640 $D=1
M424 446 750 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=33010 $D=1
M425 447 751 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=37640 $D=1
M426 444 440 446 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=33010 $D=1
M427 445 441 447 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=37640 $D=1
M428 446 78 244 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=33010 $D=1
M429 447 78 245 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=37640 $D=1
M430 248 79 446 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=33010 $D=1
M431 249 79 447 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=37640 $D=1
M432 448 79 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=33010 $D=1
M433 449 79 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=37640 $D=1
M434 6 80 450 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=33010 $D=1
M435 6 80 451 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=37640 $D=1
M436 452 81 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=33010 $D=1
M437 453 81 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=37640 $D=1
M438 454 80 234 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=33010 $D=1
M439 455 80 235 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=37640 $D=1
M440 6 454 752 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=33010 $D=1
M441 6 455 753 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=37640 $D=1
M442 456 752 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=33010 $D=1
M443 457 753 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=37640 $D=1
M444 454 450 456 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=33010 $D=1
M445 455 451 457 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=37640 $D=1
M446 456 81 244 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=33010 $D=1
M447 457 81 245 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=37640 $D=1
M448 248 82 456 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=33010 $D=1
M449 249 82 457 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=37640 $D=1
M450 458 82 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=33010 $D=1
M451 459 82 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=37640 $D=1
M452 6 83 460 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=33010 $D=1
M453 6 83 461 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=37640 $D=1
M454 462 84 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=33010 $D=1
M455 463 84 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=37640 $D=1
M456 464 83 234 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=33010 $D=1
M457 465 83 235 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=37640 $D=1
M458 6 464 754 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=33010 $D=1
M459 6 465 755 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=37640 $D=1
M460 466 754 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=33010 $D=1
M461 467 755 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=37640 $D=1
M462 464 460 466 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=33010 $D=1
M463 465 461 467 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=37640 $D=1
M464 466 84 244 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=33010 $D=1
M465 467 84 245 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=37640 $D=1
M466 248 85 466 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=33010 $D=1
M467 249 85 467 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=37640 $D=1
M468 468 85 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=33010 $D=1
M469 469 85 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=37640 $D=1
M470 6 86 470 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=33010 $D=1
M471 6 86 471 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=37640 $D=1
M472 472 87 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=33010 $D=1
M473 473 87 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=37640 $D=1
M474 474 86 234 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=33010 $D=1
M475 475 86 235 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=37640 $D=1
M476 6 474 756 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=33010 $D=1
M477 6 475 757 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=37640 $D=1
M478 476 756 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=33010 $D=1
M479 477 757 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=37640 $D=1
M480 474 470 476 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=33010 $D=1
M481 475 471 477 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=37640 $D=1
M482 476 87 244 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=33010 $D=1
M483 477 87 245 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=37640 $D=1
M484 248 88 476 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=33010 $D=1
M485 249 88 477 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=37640 $D=1
M486 478 88 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=33010 $D=1
M487 479 88 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=37640 $D=1
M488 6 89 480 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=33010 $D=1
M489 6 89 481 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=37640 $D=1
M490 482 90 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=33010 $D=1
M491 483 90 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=37640 $D=1
M492 484 89 234 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=33010 $D=1
M493 485 89 235 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=37640 $D=1
M494 6 484 758 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=33010 $D=1
M495 6 485 759 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=37640 $D=1
M496 486 758 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=33010 $D=1
M497 487 759 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=37640 $D=1
M498 484 480 486 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=33010 $D=1
M499 485 481 487 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=37640 $D=1
M500 486 90 244 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=33010 $D=1
M501 487 90 245 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=37640 $D=1
M502 248 91 486 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=33010 $D=1
M503 249 91 487 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=37640 $D=1
M504 488 91 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=33010 $D=1
M505 489 91 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=37640 $D=1
M506 6 92 490 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=33010 $D=1
M507 6 92 491 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=37640 $D=1
M508 492 93 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=33010 $D=1
M509 493 93 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=37640 $D=1
M510 494 92 234 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=33010 $D=1
M511 495 92 235 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=37640 $D=1
M512 6 494 760 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=33010 $D=1
M513 6 495 761 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=37640 $D=1
M514 496 760 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=33010 $D=1
M515 497 761 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=37640 $D=1
M516 494 490 496 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=33010 $D=1
M517 495 491 497 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=37640 $D=1
M518 496 93 244 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=33010 $D=1
M519 497 93 245 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=37640 $D=1
M520 248 94 496 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=33010 $D=1
M521 249 94 497 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=37640 $D=1
M522 498 94 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=33010 $D=1
M523 499 94 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=37640 $D=1
M524 6 95 500 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=33010 $D=1
M525 6 95 501 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=37640 $D=1
M526 502 96 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=33010 $D=1
M527 503 96 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=37640 $D=1
M528 504 95 234 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=33010 $D=1
M529 505 95 235 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=37640 $D=1
M530 6 504 762 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=33010 $D=1
M531 6 505 763 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=37640 $D=1
M532 506 762 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=33010 $D=1
M533 507 763 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=37640 $D=1
M534 504 500 506 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=33010 $D=1
M535 505 501 507 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=37640 $D=1
M536 506 96 244 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=33010 $D=1
M537 507 96 245 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=37640 $D=1
M538 248 97 506 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=33010 $D=1
M539 249 97 507 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=37640 $D=1
M540 508 97 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=33010 $D=1
M541 509 97 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=37640 $D=1
M542 6 98 510 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=33010 $D=1
M543 6 98 511 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=37640 $D=1
M544 512 99 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=33010 $D=1
M545 513 99 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=37640 $D=1
M546 514 98 234 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=33010 $D=1
M547 515 98 235 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=37640 $D=1
M548 6 514 764 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=33010 $D=1
M549 6 515 765 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=37640 $D=1
M550 516 764 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=33010 $D=1
M551 517 765 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=37640 $D=1
M552 514 510 516 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=33010 $D=1
M553 515 511 517 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=37640 $D=1
M554 516 99 244 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=33010 $D=1
M555 517 99 245 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=37640 $D=1
M556 248 100 516 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=33010 $D=1
M557 249 100 517 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=37640 $D=1
M558 518 100 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=33010 $D=1
M559 519 100 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=37640 $D=1
M560 6 101 520 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=33010 $D=1
M561 6 101 521 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=37640 $D=1
M562 522 102 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=33010 $D=1
M563 523 102 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=37640 $D=1
M564 524 101 234 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=33010 $D=1
M565 525 101 235 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=37640 $D=1
M566 6 524 766 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=33010 $D=1
M567 6 525 767 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=37640 $D=1
M568 526 766 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=33010 $D=1
M569 527 767 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=37640 $D=1
M570 524 520 526 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=33010 $D=1
M571 525 521 527 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=37640 $D=1
M572 526 102 244 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=33010 $D=1
M573 527 102 245 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=37640 $D=1
M574 248 103 526 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=33010 $D=1
M575 249 103 527 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=37640 $D=1
M576 528 103 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=33010 $D=1
M577 529 103 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=37640 $D=1
M578 6 104 530 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=33010 $D=1
M579 6 104 531 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=37640 $D=1
M580 532 105 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=33010 $D=1
M581 533 105 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=37640 $D=1
M582 534 104 234 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=33010 $D=1
M583 535 104 235 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=37640 $D=1
M584 6 534 768 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=33010 $D=1
M585 6 535 769 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=37640 $D=1
M586 536 768 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=33010 $D=1
M587 537 769 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=37640 $D=1
M588 534 530 536 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=33010 $D=1
M589 535 531 537 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=37640 $D=1
M590 536 105 244 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=33010 $D=1
M591 537 105 245 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=37640 $D=1
M592 248 109 536 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=33010 $D=1
M593 249 109 537 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=37640 $D=1
M594 538 109 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=33010 $D=1
M595 539 109 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=37640 $D=1
M596 6 111 540 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=33010 $D=1
M597 6 111 541 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=37640 $D=1
M598 542 112 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=33010 $D=1
M599 543 112 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=37640 $D=1
M600 544 111 234 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=33010 $D=1
M601 545 111 235 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=37640 $D=1
M602 6 544 770 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=33010 $D=1
M603 6 545 771 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=37640 $D=1
M604 546 770 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=33010 $D=1
M605 547 771 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=37640 $D=1
M606 544 540 546 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=33010 $D=1
M607 545 541 547 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=37640 $D=1
M608 546 112 244 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=33010 $D=1
M609 547 112 245 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=37640 $D=1
M610 248 115 546 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=33010 $D=1
M611 249 115 547 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=37640 $D=1
M612 548 115 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=33010 $D=1
M613 549 115 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=37640 $D=1
M614 6 116 550 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=33010 $D=1
M615 6 116 551 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=37640 $D=1
M616 552 117 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=33010 $D=1
M617 553 117 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=37640 $D=1
M618 6 117 244 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=33010 $D=1
M619 6 117 245 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=37640 $D=1
M620 248 116 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=33010 $D=1
M621 249 116 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=37640 $D=1
M622 6 556 554 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=33010 $D=1
M623 6 557 555 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=37640 $D=1
M624 556 118 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=33010 $D=1
M625 557 118 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=37640 $D=1
M626 772 244 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=33010 $D=1
M627 773 245 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=37640 $D=1
M628 558 554 772 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=33010 $D=1
M629 559 555 773 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=37640 $D=1
M630 6 558 560 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=33010 $D=1
M631 6 559 561 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=37640 $D=1
M632 774 560 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=33010 $D=1
M633 775 561 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=37640 $D=1
M634 558 556 774 6 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=33010 $D=1
M635 559 557 775 6 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=37640 $D=1
M636 6 564 562 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=33010 $D=1
M637 6 565 563 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=37640 $D=1
M638 564 118 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=33010 $D=1
M639 565 118 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=37640 $D=1
M640 776 248 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=33010 $D=1
M641 777 249 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=37640 $D=1
M642 566 562 776 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=33010 $D=1
M643 567 563 777 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=37640 $D=1
M644 6 566 119 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=33010 $D=1
M645 6 567 120 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=37640 $D=1
M646 778 119 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=33010 $D=1
M647 779 120 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=37640 $D=1
M648 566 564 778 6 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=33010 $D=1
M649 567 565 779 6 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=37640 $D=1
M650 568 121 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=33010 $D=1
M651 569 121 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=37640 $D=1
M652 570 568 560 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=33010 $D=1
M653 571 569 561 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=37640 $D=1
M654 122 121 570 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=33010 $D=1
M655 123 121 571 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=37640 $D=1
M656 572 124 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=33010 $D=1
M657 573 124 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=37640 $D=1
M658 574 572 119 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=33010 $D=1
M659 575 573 120 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=37640 $D=1
M660 780 124 574 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=33010 $D=1
M661 781 124 575 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=37640 $D=1
M662 6 119 780 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=33010 $D=1
M663 6 120 781 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=37640 $D=1
M664 576 125 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=33010 $D=1
M665 577 125 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=37640 $D=1
M666 578 576 574 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=33010 $D=1
M667 579 577 575 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=37640 $D=1
M668 11 125 578 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=33010 $D=1
M669 12 125 579 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=37640 $D=1
M670 581 580 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=33010 $D=1
M671 582 126 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=37640 $D=1
M672 6 585 583 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=33010 $D=1
M673 6 586 584 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=37640 $D=1
M674 587 570 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=33010 $D=1
M675 588 571 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=37640 $D=1
M676 585 587 580 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=33010 $D=1
M677 586 588 126 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=37640 $D=1
M678 581 570 585 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=33010 $D=1
M679 582 571 586 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=37640 $D=1
M680 589 583 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=33010 $D=1
M681 590 584 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=37640 $D=1
M682 127 589 578 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=33010 $D=1
M683 580 590 579 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=37640 $D=1
M684 570 583 127 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=33010 $D=1
M685 571 584 580 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=37640 $D=1
M686 591 127 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=33010 $D=1
M687 592 580 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=37640 $D=1
M688 593 583 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=33010 $D=1
M689 594 584 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=37640 $D=1
M690 595 593 591 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=33010 $D=1
M691 596 594 592 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=37640 $D=1
M692 578 583 595 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=33010 $D=1
M693 579 584 596 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=37640 $D=1
M694 597 570 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=33010 $D=1
M695 598 571 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=37640 $D=1
M696 6 578 597 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=33010 $D=1
M697 6 579 598 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=37640 $D=1
M698 599 595 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=33010 $D=1
M699 600 596 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=37640 $D=1
M700 800 570 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=33010 $D=1
M701 801 571 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=37640 $D=1
M702 601 578 800 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=33010 $D=1
M703 602 579 801 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=37640 $D=1
M704 802 570 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=33010 $D=1
M705 803 571 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=37640 $D=1
M706 603 578 802 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=33010 $D=1
M707 604 579 803 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=37640 $D=1
M708 607 570 605 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=33010 $D=1
M709 608 571 606 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=37640 $D=1
M710 605 578 607 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=33010 $D=1
M711 606 579 608 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=37640 $D=1
M712 6 603 605 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=33010 $D=1
M713 6 604 606 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=37640 $D=1
M714 609 130 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=33010 $D=1
M715 610 130 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=37640 $D=1
M716 611 609 597 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=33010 $D=1
M717 612 610 598 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=37640 $D=1
M718 601 130 611 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=33010 $D=1
M719 602 130 612 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=37640 $D=1
M720 613 609 599 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=33010 $D=1
M721 614 610 600 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=37640 $D=1
M722 607 130 613 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=33010 $D=1
M723 608 130 614 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=37640 $D=1
M724 615 131 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=33010 $D=1
M725 616 131 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=37640 $D=1
M726 617 615 613 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=33010 $D=1
M727 618 616 614 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=37640 $D=1
M728 611 131 617 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=33010 $D=1
M729 612 131 618 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=37640 $D=1
M730 13 617 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=33010 $D=1
M731 14 618 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=37640 $D=1
M732 619 132 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=33010 $D=1
M733 620 132 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=37640 $D=1
M734 621 619 133 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=33010 $D=1
M735 622 620 134 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=37640 $D=1
M736 135 132 621 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=33010 $D=1
M737 136 132 622 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=37640 $D=1
M738 623 132 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=33010 $D=1
M739 624 132 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=37640 $D=1
M740 625 623 137 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=33010 $D=1
M741 626 624 138 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=37640 $D=1
M742 139 132 625 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=33010 $D=1
M743 140 132 626 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=37640 $D=1
M744 627 132 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=33010 $D=1
M745 628 132 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=37640 $D=1
M746 629 627 128 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=33010 $D=1
M747 630 628 129 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=37640 $D=1
M748 141 132 629 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=33010 $D=1
M749 108 132 630 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=37640 $D=1
M750 631 132 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=33010 $D=1
M751 632 132 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=37640 $D=1
M752 633 631 142 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=33010 $D=1
M753 634 632 143 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=37640 $D=1
M754 144 132 633 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=33010 $D=1
M755 145 132 634 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=37640 $D=1
M756 635 132 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=33010 $D=1
M757 636 132 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=37640 $D=1
M758 637 635 146 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=33010 $D=1
M759 638 636 147 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=37640 $D=1
M760 144 132 637 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=33010 $D=1
M761 144 132 638 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=37640 $D=1
M762 6 570 782 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=33010 $D=1
M763 6 571 783 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=37640 $D=1
M764 136 782 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=33010 $D=1
M765 133 783 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=37640 $D=1
M766 639 148 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=33010 $D=1
M767 640 148 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=37640 $D=1
M768 149 639 136 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=33010 $D=1
M769 150 640 133 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=37640 $D=1
M770 621 148 149 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=33010 $D=1
M771 622 148 150 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=37640 $D=1
M772 641 151 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=33010 $D=1
M773 642 151 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=37640 $D=1
M774 152 641 149 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=33010 $D=1
M775 113 642 150 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=37640 $D=1
M776 625 151 152 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=33010 $D=1
M777 626 151 113 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=37640 $D=1
M778 643 153 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=33010 $D=1
M779 644 153 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=37640 $D=1
M780 154 643 152 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=33010 $D=1
M781 106 644 113 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=37640 $D=1
M782 629 153 154 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=33010 $D=1
M783 630 153 106 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=37640 $D=1
M784 645 155 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=33010 $D=1
M785 646 155 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=37640 $D=1
M786 156 645 154 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=33010 $D=1
M787 157 646 106 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=37640 $D=1
M788 633 155 156 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=33010 $D=1
M789 634 155 157 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=37640 $D=1
M790 647 158 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=33010 $D=1
M791 648 158 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=37640 $D=1
M792 220 647 156 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=33010 $D=1
M793 221 648 157 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=37640 $D=1
M794 637 158 220 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=33010 $D=1
M795 638 158 221 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=37640 $D=1
M796 649 159 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=33010 $D=1
M797 650 159 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=37640 $D=1
M798 651 649 119 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=33010 $D=1
M799 652 650 120 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=37640 $D=1
M800 11 159 651 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=33010 $D=1
M801 12 159 652 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=37640 $D=1
M802 804 560 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=33010 $D=1
M803 805 561 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=37640 $D=1
M804 653 651 804 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=33010 $D=1
M805 654 652 805 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=37640 $D=1
M806 657 560 655 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=33010 $D=1
M807 658 561 656 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=37640 $D=1
M808 655 651 657 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=33010 $D=1
M809 656 652 658 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=37640 $D=1
M810 6 653 655 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=33010 $D=1
M811 6 654 656 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=37640 $D=1
M812 806 160 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=33010 $D=1
M813 807 659 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=37640 $D=1
M814 784 657 806 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=33010 $D=1
M815 785 658 807 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=37640 $D=1
M816 659 784 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=33010 $D=1
M817 161 785 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=37640 $D=1
M818 660 560 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=33010 $D=1
M819 661 561 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=37640 $D=1
M820 6 662 660 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=33010 $D=1
M821 6 663 661 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=37640 $D=1
M822 662 651 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=33010 $D=1
M823 663 652 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=37640 $D=1
M824 808 660 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=33010 $D=1
M825 809 661 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=37640 $D=1
M826 664 160 808 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=33010 $D=1
M827 665 659 809 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=37640 $D=1
M828 667 162 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=33010 $D=1
M829 668 666 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=37640 $D=1
M830 810 664 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=33010 $D=1
M831 811 665 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=37640 $D=1
M832 666 667 810 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=33010 $D=1
M833 163 668 811 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=37640 $D=1
M834 670 669 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=33010 $D=1
M835 671 164 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=37640 $D=1
M836 6 674 672 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=33010 $D=1
M837 6 675 673 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=37640 $D=1
M838 676 122 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=33010 $D=1
M839 677 123 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=37640 $D=1
M840 674 676 669 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=33010 $D=1
M841 675 677 164 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=37640 $D=1
M842 670 122 674 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=33010 $D=1
M843 671 123 675 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=37640 $D=1
M844 678 672 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=33010 $D=1
M845 679 673 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=37640 $D=1
M846 165 678 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=33010 $D=1
M847 669 679 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=37640 $D=1
M848 122 672 165 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=33010 $D=1
M849 123 673 669 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=37640 $D=1
M850 680 165 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=33010 $D=1
M851 681 669 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=37640 $D=1
M852 682 672 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=33010 $D=1
M853 683 673 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=37640 $D=1
M854 222 682 680 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=33010 $D=1
M855 223 683 681 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=37640 $D=1
M856 6 672 222 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=33010 $D=1
M857 6 673 223 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=37640 $D=1
M858 684 166 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=33010 $D=1
M859 685 166 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=37640 $D=1
M860 686 684 222 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=33010 $D=1
M861 687 685 223 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=37640 $D=1
M862 13 166 686 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=33010 $D=1
M863 14 166 687 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=37640 $D=1
M864 688 167 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=33010 $D=1
M865 689 167 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=37640 $D=1
M866 690 688 686 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=33010 $D=1
M867 691 689 687 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=37640 $D=1
M868 6 167 690 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=33010 $D=1
M869 6 167 691 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=37640 $D=1
M870 692 118 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=33010 $D=1
M871 693 118 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=37640 $D=1
M872 6 692 694 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=33010 $D=1
M873 6 693 695 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=37640 $D=1
M874 696 118 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=33010 $D=1
M875 697 118 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=37640 $D=1
M876 698 692 690 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=33010 $D=1
M877 699 693 691 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=37640 $D=1
M878 6 698 786 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=33010 $D=1
M879 6 699 787 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=37640 $D=1
M880 700 786 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=33010 $D=1
M881 701 787 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=37640 $D=1
M882 698 694 700 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=33010 $D=1
M883 699 695 701 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=37640 $D=1
M884 702 118 700 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=33010 $D=1
M885 703 118 701 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=37640 $D=1
M886 6 706 704 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=33010 $D=1
M887 6 707 705 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=37640 $D=1
M888 706 118 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=33010 $D=1
M889 707 118 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=37640 $D=1
M890 788 702 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=33010 $D=1
M891 789 703 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=37640 $D=1
M892 708 704 788 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=33010 $D=1
M893 709 705 789 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=37640 $D=1
M894 6 708 122 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=33010 $D=1
M895 6 709 123 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=37640 $D=1
M896 790 122 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=33010 $D=1
M897 791 123 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=37640 $D=1
M898 708 706 790 6 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=33010 $D=1
M899 709 707 791 6 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=37640 $D=1
M900 196 1 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=34260 $D=0
M901 197 1 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=38890 $D=0
M902 198 1 2 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=34260 $D=0
M903 199 1 3 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=38890 $D=0
M904 6 196 198 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=34260 $D=0
M905 6 197 199 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=38890 $D=0
M906 200 1 4 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=34260 $D=0
M907 201 1 4 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=38890 $D=0
M908 5 196 200 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=34260 $D=0
M909 5 197 201 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=38890 $D=0
M910 202 1 6 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=34260 $D=0
M911 203 1 6 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=38890 $D=0
M912 6 196 202 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=34260 $D=0
M913 6 197 203 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=38890 $D=0
M914 206 7 202 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=34260 $D=0
M915 207 7 203 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=38890 $D=0
M916 204 7 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=34260 $D=0
M917 205 7 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=38890 $D=0
M918 208 7 200 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=34260 $D=0
M919 209 7 201 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=38890 $D=0
M920 198 204 208 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=34260 $D=0
M921 199 205 209 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=38890 $D=0
M922 210 8 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=34260 $D=0
M923 211 8 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=38890 $D=0
M924 212 8 208 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=34260 $D=0
M925 213 8 209 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=38890 $D=0
M926 206 210 212 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=34260 $D=0
M927 207 211 213 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=38890 $D=0
M928 214 10 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=34260 $D=0
M929 215 10 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=38890 $D=0
M930 216 10 6 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=34260 $D=0
M931 217 10 6 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=38890 $D=0
M932 11 214 216 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=34260 $D=0
M933 12 215 217 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=38890 $D=0
M934 218 10 13 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=34260 $D=0
M935 219 10 14 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=38890 $D=0
M936 220 214 218 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=34260 $D=0
M937 221 215 219 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=38890 $D=0
M938 224 10 222 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=34260 $D=0
M939 225 10 223 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=38890 $D=0
M940 212 214 224 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=34260 $D=0
M941 213 215 225 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=38890 $D=0
M942 228 15 224 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=34260 $D=0
M943 229 15 225 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=38890 $D=0
M944 226 15 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=34260 $D=0
M945 227 15 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=38890 $D=0
M946 230 15 218 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=34260 $D=0
M947 231 15 219 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=38890 $D=0
M948 216 226 230 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=34260 $D=0
M949 217 227 231 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=38890 $D=0
M950 232 16 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=34260 $D=0
M951 233 16 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=38890 $D=0
M952 234 16 230 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=34260 $D=0
M953 235 16 231 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=38890 $D=0
M954 228 232 234 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=34260 $D=0
M955 229 233 235 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=38890 $D=0
M956 9 17 236 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=34260 $D=0
M957 9 17 237 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=38890 $D=0
M958 238 18 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=34260 $D=0
M959 239 18 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=38890 $D=0
M960 240 236 234 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=34260 $D=0
M961 241 237 235 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=38890 $D=0
M962 9 240 710 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=34260 $D=0
M963 9 241 711 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=38890 $D=0
M964 242 710 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=34260 $D=0
M965 243 711 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=38890 $D=0
M966 240 17 242 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=34260 $D=0
M967 241 17 243 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=38890 $D=0
M968 242 238 244 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=34260 $D=0
M969 243 239 245 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=38890 $D=0
M970 248 246 242 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=34260 $D=0
M971 249 247 243 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=38890 $D=0
M972 246 19 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=34260 $D=0
M973 247 19 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=38890 $D=0
M974 9 20 250 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=34260 $D=0
M975 9 20 251 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=38890 $D=0
M976 252 21 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=34260 $D=0
M977 253 21 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=38890 $D=0
M978 254 250 234 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=34260 $D=0
M979 255 251 235 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=38890 $D=0
M980 9 254 712 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=34260 $D=0
M981 9 255 713 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=38890 $D=0
M982 256 712 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=34260 $D=0
M983 257 713 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=38890 $D=0
M984 254 20 256 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=34260 $D=0
M985 255 20 257 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=38890 $D=0
M986 256 252 244 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=34260 $D=0
M987 257 253 245 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=38890 $D=0
M988 248 258 256 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=34260 $D=0
M989 249 259 257 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=38890 $D=0
M990 258 22 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=34260 $D=0
M991 259 22 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=38890 $D=0
M992 9 23 260 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=34260 $D=0
M993 9 23 261 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=38890 $D=0
M994 262 24 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=34260 $D=0
M995 263 24 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=38890 $D=0
M996 264 260 234 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=34260 $D=0
M997 265 261 235 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=38890 $D=0
M998 9 264 714 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=34260 $D=0
M999 9 265 715 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=38890 $D=0
M1000 266 714 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=34260 $D=0
M1001 267 715 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=38890 $D=0
M1002 264 23 266 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=34260 $D=0
M1003 265 23 267 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=38890 $D=0
M1004 266 262 244 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=34260 $D=0
M1005 267 263 245 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=38890 $D=0
M1006 248 268 266 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=34260 $D=0
M1007 249 269 267 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=38890 $D=0
M1008 268 25 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=34260 $D=0
M1009 269 25 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=38890 $D=0
M1010 9 26 270 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=34260 $D=0
M1011 9 26 271 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=38890 $D=0
M1012 272 27 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=34260 $D=0
M1013 273 27 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=38890 $D=0
M1014 274 270 234 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=34260 $D=0
M1015 275 271 235 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=38890 $D=0
M1016 9 274 716 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=34260 $D=0
M1017 9 275 717 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=38890 $D=0
M1018 276 716 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=34260 $D=0
M1019 277 717 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=38890 $D=0
M1020 274 26 276 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=34260 $D=0
M1021 275 26 277 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=38890 $D=0
M1022 276 272 244 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=34260 $D=0
M1023 277 273 245 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=38890 $D=0
M1024 248 278 276 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=34260 $D=0
M1025 249 279 277 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=38890 $D=0
M1026 278 28 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=34260 $D=0
M1027 279 28 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=38890 $D=0
M1028 9 29 280 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=34260 $D=0
M1029 9 29 281 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=38890 $D=0
M1030 282 30 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=34260 $D=0
M1031 283 30 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=38890 $D=0
M1032 284 280 234 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=34260 $D=0
M1033 285 281 235 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=38890 $D=0
M1034 9 284 718 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=34260 $D=0
M1035 9 285 719 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=38890 $D=0
M1036 286 718 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=34260 $D=0
M1037 287 719 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=38890 $D=0
M1038 284 29 286 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=34260 $D=0
M1039 285 29 287 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=38890 $D=0
M1040 286 282 244 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=34260 $D=0
M1041 287 283 245 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=38890 $D=0
M1042 248 288 286 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=34260 $D=0
M1043 249 289 287 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=38890 $D=0
M1044 288 31 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=34260 $D=0
M1045 289 31 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=38890 $D=0
M1046 9 32 290 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=34260 $D=0
M1047 9 32 291 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=38890 $D=0
M1048 292 33 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=34260 $D=0
M1049 293 33 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=38890 $D=0
M1050 294 290 234 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=34260 $D=0
M1051 295 291 235 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=38890 $D=0
M1052 9 294 720 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=34260 $D=0
M1053 9 295 721 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=38890 $D=0
M1054 296 720 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=34260 $D=0
M1055 297 721 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=38890 $D=0
M1056 294 32 296 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=34260 $D=0
M1057 295 32 297 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=38890 $D=0
M1058 296 292 244 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=34260 $D=0
M1059 297 293 245 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=38890 $D=0
M1060 248 298 296 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=34260 $D=0
M1061 249 299 297 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=38890 $D=0
M1062 298 34 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=34260 $D=0
M1063 299 34 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=38890 $D=0
M1064 9 35 300 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=34260 $D=0
M1065 9 35 301 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=38890 $D=0
M1066 302 36 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=34260 $D=0
M1067 303 36 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=38890 $D=0
M1068 304 300 234 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=34260 $D=0
M1069 305 301 235 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=38890 $D=0
M1070 9 304 722 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=34260 $D=0
M1071 9 305 723 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=38890 $D=0
M1072 306 722 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=34260 $D=0
M1073 307 723 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=38890 $D=0
M1074 304 35 306 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=34260 $D=0
M1075 305 35 307 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=38890 $D=0
M1076 306 302 244 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=34260 $D=0
M1077 307 303 245 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=38890 $D=0
M1078 248 308 306 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=34260 $D=0
M1079 249 309 307 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=38890 $D=0
M1080 308 37 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=34260 $D=0
M1081 309 37 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=38890 $D=0
M1082 9 38 310 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=34260 $D=0
M1083 9 38 311 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=38890 $D=0
M1084 312 39 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=34260 $D=0
M1085 313 39 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=38890 $D=0
M1086 314 310 234 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=34260 $D=0
M1087 315 311 235 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=38890 $D=0
M1088 9 314 724 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=34260 $D=0
M1089 9 315 725 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=38890 $D=0
M1090 316 724 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=34260 $D=0
M1091 317 725 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=38890 $D=0
M1092 314 38 316 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=34260 $D=0
M1093 315 38 317 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=38890 $D=0
M1094 316 312 244 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=34260 $D=0
M1095 317 313 245 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=38890 $D=0
M1096 248 318 316 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=34260 $D=0
M1097 249 319 317 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=38890 $D=0
M1098 318 40 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=34260 $D=0
M1099 319 40 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=38890 $D=0
M1100 9 41 320 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=34260 $D=0
M1101 9 41 321 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=38890 $D=0
M1102 322 42 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=34260 $D=0
M1103 323 42 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=38890 $D=0
M1104 324 320 234 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=34260 $D=0
M1105 325 321 235 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=38890 $D=0
M1106 9 324 726 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=34260 $D=0
M1107 9 325 727 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=38890 $D=0
M1108 326 726 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=34260 $D=0
M1109 327 727 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=38890 $D=0
M1110 324 41 326 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=34260 $D=0
M1111 325 41 327 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=38890 $D=0
M1112 326 322 244 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=34260 $D=0
M1113 327 323 245 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=38890 $D=0
M1114 248 328 326 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=34260 $D=0
M1115 249 329 327 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=38890 $D=0
M1116 328 43 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=34260 $D=0
M1117 329 43 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=38890 $D=0
M1118 9 44 330 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=34260 $D=0
M1119 9 44 331 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=38890 $D=0
M1120 332 45 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=34260 $D=0
M1121 333 45 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=38890 $D=0
M1122 334 330 234 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=34260 $D=0
M1123 335 331 235 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=38890 $D=0
M1124 9 334 728 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=34260 $D=0
M1125 9 335 729 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=38890 $D=0
M1126 336 728 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=34260 $D=0
M1127 337 729 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=38890 $D=0
M1128 334 44 336 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=34260 $D=0
M1129 335 44 337 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=38890 $D=0
M1130 336 332 244 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=34260 $D=0
M1131 337 333 245 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=38890 $D=0
M1132 248 338 336 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=34260 $D=0
M1133 249 339 337 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=38890 $D=0
M1134 338 46 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=34260 $D=0
M1135 339 46 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=38890 $D=0
M1136 9 47 340 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=34260 $D=0
M1137 9 47 341 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=38890 $D=0
M1138 342 48 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=34260 $D=0
M1139 343 48 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=38890 $D=0
M1140 344 340 234 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=34260 $D=0
M1141 345 341 235 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=38890 $D=0
M1142 9 344 730 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=34260 $D=0
M1143 9 345 731 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=38890 $D=0
M1144 346 730 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=34260 $D=0
M1145 347 731 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=38890 $D=0
M1146 344 47 346 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=34260 $D=0
M1147 345 47 347 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=38890 $D=0
M1148 346 342 244 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=34260 $D=0
M1149 347 343 245 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=38890 $D=0
M1150 248 348 346 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=34260 $D=0
M1151 249 349 347 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=38890 $D=0
M1152 348 49 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=34260 $D=0
M1153 349 49 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=38890 $D=0
M1154 9 50 350 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=34260 $D=0
M1155 9 50 351 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=38890 $D=0
M1156 352 51 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=34260 $D=0
M1157 353 51 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=38890 $D=0
M1158 354 350 234 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=34260 $D=0
M1159 355 351 235 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=38890 $D=0
M1160 9 354 732 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=34260 $D=0
M1161 9 355 733 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=38890 $D=0
M1162 356 732 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=34260 $D=0
M1163 357 733 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=38890 $D=0
M1164 354 50 356 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=34260 $D=0
M1165 355 50 357 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=38890 $D=0
M1166 356 352 244 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=34260 $D=0
M1167 357 353 245 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=38890 $D=0
M1168 248 358 356 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=34260 $D=0
M1169 249 359 357 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=38890 $D=0
M1170 358 52 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=34260 $D=0
M1171 359 52 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=38890 $D=0
M1172 9 53 360 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=34260 $D=0
M1173 9 53 361 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=38890 $D=0
M1174 362 54 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=34260 $D=0
M1175 363 54 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=38890 $D=0
M1176 364 360 234 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=34260 $D=0
M1177 365 361 235 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=38890 $D=0
M1178 9 364 734 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=34260 $D=0
M1179 9 365 735 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=38890 $D=0
M1180 366 734 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=34260 $D=0
M1181 367 735 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=38890 $D=0
M1182 364 53 366 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=34260 $D=0
M1183 365 53 367 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=38890 $D=0
M1184 366 362 244 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=34260 $D=0
M1185 367 363 245 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=38890 $D=0
M1186 248 368 366 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=34260 $D=0
M1187 249 369 367 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=38890 $D=0
M1188 368 55 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=34260 $D=0
M1189 369 55 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=38890 $D=0
M1190 9 56 370 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=34260 $D=0
M1191 9 56 371 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=38890 $D=0
M1192 372 57 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=34260 $D=0
M1193 373 57 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=38890 $D=0
M1194 374 370 234 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=34260 $D=0
M1195 375 371 235 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=38890 $D=0
M1196 9 374 736 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=34260 $D=0
M1197 9 375 737 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=38890 $D=0
M1198 376 736 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=34260 $D=0
M1199 377 737 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=38890 $D=0
M1200 374 56 376 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=34260 $D=0
M1201 375 56 377 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=38890 $D=0
M1202 376 372 244 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=34260 $D=0
M1203 377 373 245 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=38890 $D=0
M1204 248 378 376 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=34260 $D=0
M1205 249 379 377 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=38890 $D=0
M1206 378 58 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=34260 $D=0
M1207 379 58 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=38890 $D=0
M1208 9 59 380 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=34260 $D=0
M1209 9 59 381 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=38890 $D=0
M1210 382 60 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=34260 $D=0
M1211 383 60 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=38890 $D=0
M1212 384 380 234 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=34260 $D=0
M1213 385 381 235 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=38890 $D=0
M1214 9 384 738 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=34260 $D=0
M1215 9 385 739 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=38890 $D=0
M1216 386 738 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=34260 $D=0
M1217 387 739 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=38890 $D=0
M1218 384 59 386 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=34260 $D=0
M1219 385 59 387 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=38890 $D=0
M1220 386 382 244 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=34260 $D=0
M1221 387 383 245 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=38890 $D=0
M1222 248 388 386 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=34260 $D=0
M1223 249 389 387 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=38890 $D=0
M1224 388 61 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=34260 $D=0
M1225 389 61 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=38890 $D=0
M1226 9 62 390 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=34260 $D=0
M1227 9 62 391 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=38890 $D=0
M1228 392 63 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=34260 $D=0
M1229 393 63 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=38890 $D=0
M1230 394 390 234 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=34260 $D=0
M1231 395 391 235 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=38890 $D=0
M1232 9 394 740 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=34260 $D=0
M1233 9 395 741 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=38890 $D=0
M1234 396 740 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=34260 $D=0
M1235 397 741 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=38890 $D=0
M1236 394 62 396 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=34260 $D=0
M1237 395 62 397 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=38890 $D=0
M1238 396 392 244 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=34260 $D=0
M1239 397 393 245 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=38890 $D=0
M1240 248 398 396 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=34260 $D=0
M1241 249 399 397 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=38890 $D=0
M1242 398 64 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=34260 $D=0
M1243 399 64 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=38890 $D=0
M1244 9 65 400 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=34260 $D=0
M1245 9 65 401 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=38890 $D=0
M1246 402 66 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=34260 $D=0
M1247 403 66 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=38890 $D=0
M1248 404 400 234 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=34260 $D=0
M1249 405 401 235 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=38890 $D=0
M1250 9 404 742 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=34260 $D=0
M1251 9 405 743 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=38890 $D=0
M1252 406 742 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=34260 $D=0
M1253 407 743 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=38890 $D=0
M1254 404 65 406 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=34260 $D=0
M1255 405 65 407 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=38890 $D=0
M1256 406 402 244 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=34260 $D=0
M1257 407 403 245 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=38890 $D=0
M1258 248 408 406 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=34260 $D=0
M1259 249 409 407 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=38890 $D=0
M1260 408 67 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=34260 $D=0
M1261 409 67 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=38890 $D=0
M1262 9 68 410 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=34260 $D=0
M1263 9 68 411 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=38890 $D=0
M1264 412 69 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=34260 $D=0
M1265 413 69 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=38890 $D=0
M1266 414 410 234 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=34260 $D=0
M1267 415 411 235 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=38890 $D=0
M1268 9 414 744 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=34260 $D=0
M1269 9 415 745 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=38890 $D=0
M1270 416 744 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=34260 $D=0
M1271 417 745 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=38890 $D=0
M1272 414 68 416 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=34260 $D=0
M1273 415 68 417 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=38890 $D=0
M1274 416 412 244 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=34260 $D=0
M1275 417 413 245 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=38890 $D=0
M1276 248 418 416 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=34260 $D=0
M1277 249 419 417 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=38890 $D=0
M1278 418 70 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=34260 $D=0
M1279 419 70 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=38890 $D=0
M1280 9 71 420 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=34260 $D=0
M1281 9 71 421 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=38890 $D=0
M1282 422 72 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=34260 $D=0
M1283 423 72 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=38890 $D=0
M1284 424 420 234 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=34260 $D=0
M1285 425 421 235 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=38890 $D=0
M1286 9 424 746 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=34260 $D=0
M1287 9 425 747 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=38890 $D=0
M1288 426 746 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=34260 $D=0
M1289 427 747 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=38890 $D=0
M1290 424 71 426 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=34260 $D=0
M1291 425 71 427 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=38890 $D=0
M1292 426 422 244 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=34260 $D=0
M1293 427 423 245 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=38890 $D=0
M1294 248 428 426 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=34260 $D=0
M1295 249 429 427 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=38890 $D=0
M1296 428 73 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=34260 $D=0
M1297 429 73 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=38890 $D=0
M1298 9 74 430 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=34260 $D=0
M1299 9 74 431 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=38890 $D=0
M1300 432 75 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=34260 $D=0
M1301 433 75 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=38890 $D=0
M1302 434 430 234 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=34260 $D=0
M1303 435 431 235 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=38890 $D=0
M1304 9 434 748 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=34260 $D=0
M1305 9 435 749 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=38890 $D=0
M1306 436 748 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=34260 $D=0
M1307 437 749 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=38890 $D=0
M1308 434 74 436 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=34260 $D=0
M1309 435 74 437 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=38890 $D=0
M1310 436 432 244 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=34260 $D=0
M1311 437 433 245 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=38890 $D=0
M1312 248 438 436 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=34260 $D=0
M1313 249 439 437 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=38890 $D=0
M1314 438 76 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=34260 $D=0
M1315 439 76 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=38890 $D=0
M1316 9 77 440 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=34260 $D=0
M1317 9 77 441 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=38890 $D=0
M1318 442 78 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=34260 $D=0
M1319 443 78 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=38890 $D=0
M1320 444 440 234 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=34260 $D=0
M1321 445 441 235 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=38890 $D=0
M1322 9 444 750 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=34260 $D=0
M1323 9 445 751 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=38890 $D=0
M1324 446 750 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=34260 $D=0
M1325 447 751 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=38890 $D=0
M1326 444 77 446 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=34260 $D=0
M1327 445 77 447 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=38890 $D=0
M1328 446 442 244 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=34260 $D=0
M1329 447 443 245 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=38890 $D=0
M1330 248 448 446 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=34260 $D=0
M1331 249 449 447 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=38890 $D=0
M1332 448 79 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=34260 $D=0
M1333 449 79 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=38890 $D=0
M1334 9 80 450 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=34260 $D=0
M1335 9 80 451 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=38890 $D=0
M1336 452 81 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=34260 $D=0
M1337 453 81 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=38890 $D=0
M1338 454 450 234 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=34260 $D=0
M1339 455 451 235 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=38890 $D=0
M1340 9 454 752 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=34260 $D=0
M1341 9 455 753 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=38890 $D=0
M1342 456 752 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=34260 $D=0
M1343 457 753 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=38890 $D=0
M1344 454 80 456 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=34260 $D=0
M1345 455 80 457 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=38890 $D=0
M1346 456 452 244 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=34260 $D=0
M1347 457 453 245 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=38890 $D=0
M1348 248 458 456 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=34260 $D=0
M1349 249 459 457 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=38890 $D=0
M1350 458 82 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=34260 $D=0
M1351 459 82 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=38890 $D=0
M1352 9 83 460 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=34260 $D=0
M1353 9 83 461 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=38890 $D=0
M1354 462 84 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=34260 $D=0
M1355 463 84 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=38890 $D=0
M1356 464 460 234 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=34260 $D=0
M1357 465 461 235 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=38890 $D=0
M1358 9 464 754 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=34260 $D=0
M1359 9 465 755 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=38890 $D=0
M1360 466 754 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=34260 $D=0
M1361 467 755 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=38890 $D=0
M1362 464 83 466 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=34260 $D=0
M1363 465 83 467 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=38890 $D=0
M1364 466 462 244 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=34260 $D=0
M1365 467 463 245 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=38890 $D=0
M1366 248 468 466 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=34260 $D=0
M1367 249 469 467 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=38890 $D=0
M1368 468 85 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=34260 $D=0
M1369 469 85 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=38890 $D=0
M1370 9 86 470 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=34260 $D=0
M1371 9 86 471 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=38890 $D=0
M1372 472 87 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=34260 $D=0
M1373 473 87 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=38890 $D=0
M1374 474 470 234 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=34260 $D=0
M1375 475 471 235 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=38890 $D=0
M1376 9 474 756 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=34260 $D=0
M1377 9 475 757 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=38890 $D=0
M1378 476 756 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=34260 $D=0
M1379 477 757 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=38890 $D=0
M1380 474 86 476 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=34260 $D=0
M1381 475 86 477 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=38890 $D=0
M1382 476 472 244 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=34260 $D=0
M1383 477 473 245 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=38890 $D=0
M1384 248 478 476 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=34260 $D=0
M1385 249 479 477 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=38890 $D=0
M1386 478 88 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=34260 $D=0
M1387 479 88 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=38890 $D=0
M1388 9 89 480 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=34260 $D=0
M1389 9 89 481 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=38890 $D=0
M1390 482 90 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=34260 $D=0
M1391 483 90 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=38890 $D=0
M1392 484 480 234 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=34260 $D=0
M1393 485 481 235 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=38890 $D=0
M1394 9 484 758 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=34260 $D=0
M1395 9 485 759 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=38890 $D=0
M1396 486 758 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=34260 $D=0
M1397 487 759 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=38890 $D=0
M1398 484 89 486 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=34260 $D=0
M1399 485 89 487 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=38890 $D=0
M1400 486 482 244 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=34260 $D=0
M1401 487 483 245 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=38890 $D=0
M1402 248 488 486 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=34260 $D=0
M1403 249 489 487 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=38890 $D=0
M1404 488 91 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=34260 $D=0
M1405 489 91 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=38890 $D=0
M1406 9 92 490 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=34260 $D=0
M1407 9 92 491 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=38890 $D=0
M1408 492 93 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=34260 $D=0
M1409 493 93 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=38890 $D=0
M1410 494 490 234 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=34260 $D=0
M1411 495 491 235 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=38890 $D=0
M1412 9 494 760 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=34260 $D=0
M1413 9 495 761 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=38890 $D=0
M1414 496 760 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=34260 $D=0
M1415 497 761 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=38890 $D=0
M1416 494 92 496 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=34260 $D=0
M1417 495 92 497 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=38890 $D=0
M1418 496 492 244 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=34260 $D=0
M1419 497 493 245 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=38890 $D=0
M1420 248 498 496 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=34260 $D=0
M1421 249 499 497 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=38890 $D=0
M1422 498 94 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=34260 $D=0
M1423 499 94 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=38890 $D=0
M1424 9 95 500 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=34260 $D=0
M1425 9 95 501 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=38890 $D=0
M1426 502 96 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=34260 $D=0
M1427 503 96 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=38890 $D=0
M1428 504 500 234 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=34260 $D=0
M1429 505 501 235 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=38890 $D=0
M1430 9 504 762 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=34260 $D=0
M1431 9 505 763 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=38890 $D=0
M1432 506 762 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=34260 $D=0
M1433 507 763 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=38890 $D=0
M1434 504 95 506 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=34260 $D=0
M1435 505 95 507 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=38890 $D=0
M1436 506 502 244 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=34260 $D=0
M1437 507 503 245 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=38890 $D=0
M1438 248 508 506 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=34260 $D=0
M1439 249 509 507 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=38890 $D=0
M1440 508 97 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=34260 $D=0
M1441 509 97 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=38890 $D=0
M1442 9 98 510 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=34260 $D=0
M1443 9 98 511 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=38890 $D=0
M1444 512 99 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=34260 $D=0
M1445 513 99 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=38890 $D=0
M1446 514 510 234 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=34260 $D=0
M1447 515 511 235 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=38890 $D=0
M1448 9 514 764 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=34260 $D=0
M1449 9 515 765 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=38890 $D=0
M1450 516 764 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=34260 $D=0
M1451 517 765 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=38890 $D=0
M1452 514 98 516 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=34260 $D=0
M1453 515 98 517 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=38890 $D=0
M1454 516 512 244 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=34260 $D=0
M1455 517 513 245 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=38890 $D=0
M1456 248 518 516 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=34260 $D=0
M1457 249 519 517 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=38890 $D=0
M1458 518 100 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=34260 $D=0
M1459 519 100 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=38890 $D=0
M1460 9 101 520 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=34260 $D=0
M1461 9 101 521 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=38890 $D=0
M1462 522 102 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=34260 $D=0
M1463 523 102 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=38890 $D=0
M1464 524 520 234 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=34260 $D=0
M1465 525 521 235 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=38890 $D=0
M1466 9 524 766 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=34260 $D=0
M1467 9 525 767 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=38890 $D=0
M1468 526 766 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=34260 $D=0
M1469 527 767 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=38890 $D=0
M1470 524 101 526 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=34260 $D=0
M1471 525 101 527 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=38890 $D=0
M1472 526 522 244 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=34260 $D=0
M1473 527 523 245 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=38890 $D=0
M1474 248 528 526 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=34260 $D=0
M1475 249 529 527 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=38890 $D=0
M1476 528 103 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=34260 $D=0
M1477 529 103 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=38890 $D=0
M1478 9 104 530 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=34260 $D=0
M1479 9 104 531 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=38890 $D=0
M1480 532 105 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=34260 $D=0
M1481 533 105 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=38890 $D=0
M1482 534 530 234 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=34260 $D=0
M1483 535 531 235 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=38890 $D=0
M1484 9 534 768 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=34260 $D=0
M1485 9 535 769 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=38890 $D=0
M1486 536 768 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=34260 $D=0
M1487 537 769 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=38890 $D=0
M1488 534 104 536 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=34260 $D=0
M1489 535 104 537 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=38890 $D=0
M1490 536 532 244 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=34260 $D=0
M1491 537 533 245 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=38890 $D=0
M1492 248 538 536 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=34260 $D=0
M1493 249 539 537 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=38890 $D=0
M1494 538 109 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=34260 $D=0
M1495 539 109 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=38890 $D=0
M1496 9 111 540 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=34260 $D=0
M1497 9 111 541 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=38890 $D=0
M1498 542 112 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=34260 $D=0
M1499 543 112 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=38890 $D=0
M1500 544 540 234 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=34260 $D=0
M1501 545 541 235 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=38890 $D=0
M1502 9 544 770 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=34260 $D=0
M1503 9 545 771 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=38890 $D=0
M1504 546 770 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=34260 $D=0
M1505 547 771 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=38890 $D=0
M1506 544 111 546 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=34260 $D=0
M1507 545 111 547 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=38890 $D=0
M1508 546 542 244 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=34260 $D=0
M1509 547 543 245 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=38890 $D=0
M1510 248 548 546 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=34260 $D=0
M1511 249 549 547 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=38890 $D=0
M1512 548 115 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=34260 $D=0
M1513 549 115 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=38890 $D=0
M1514 9 116 550 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=34260 $D=0
M1515 9 116 551 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=38890 $D=0
M1516 552 117 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=34260 $D=0
M1517 553 117 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=38890 $D=0
M1518 6 552 244 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=34260 $D=0
M1519 6 553 245 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=38890 $D=0
M1520 248 550 6 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=34260 $D=0
M1521 249 551 6 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=38890 $D=0
M1522 9 556 554 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=34260 $D=0
M1523 9 557 555 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=38890 $D=0
M1524 556 118 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=34260 $D=0
M1525 557 118 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=38890 $D=0
M1526 772 244 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=34260 $D=0
M1527 773 245 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=38890 $D=0
M1528 558 556 772 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=34260 $D=0
M1529 559 557 773 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=38890 $D=0
M1530 9 558 560 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=34260 $D=0
M1531 9 559 561 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=38890 $D=0
M1532 774 560 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=34260 $D=0
M1533 775 561 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=38890 $D=0
M1534 558 554 774 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=34260 $D=0
M1535 559 555 775 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=38890 $D=0
M1536 9 564 562 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=34260 $D=0
M1537 9 565 563 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=38890 $D=0
M1538 564 118 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=34260 $D=0
M1539 565 118 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=38890 $D=0
M1540 776 248 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=34260 $D=0
M1541 777 249 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=38890 $D=0
M1542 566 564 776 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=34260 $D=0
M1543 567 565 777 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=38890 $D=0
M1544 9 566 119 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=34260 $D=0
M1545 9 567 120 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=38890 $D=0
M1546 778 119 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=34260 $D=0
M1547 779 120 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=38890 $D=0
M1548 566 562 778 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=34260 $D=0
M1549 567 563 779 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=38890 $D=0
M1550 568 121 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=34260 $D=0
M1551 569 121 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=38890 $D=0
M1552 570 121 560 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=34260 $D=0
M1553 571 121 561 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=38890 $D=0
M1554 122 568 570 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=34260 $D=0
M1555 123 569 571 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=38890 $D=0
M1556 572 124 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=34260 $D=0
M1557 573 124 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=38890 $D=0
M1558 574 124 119 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=34260 $D=0
M1559 575 124 120 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=38890 $D=0
M1560 780 572 574 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=34260 $D=0
M1561 781 573 575 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=38890 $D=0
M1562 9 119 780 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=34260 $D=0
M1563 9 120 781 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=38890 $D=0
M1564 576 125 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=34260 $D=0
M1565 577 125 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=38890 $D=0
M1566 578 125 574 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=34260 $D=0
M1567 579 125 575 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=38890 $D=0
M1568 11 576 578 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=34260 $D=0
M1569 12 577 579 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=38890 $D=0
M1570 581 580 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=34260 $D=0
M1571 582 126 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=38890 $D=0
M1572 9 585 583 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=34260 $D=0
M1573 9 586 584 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=38890 $D=0
M1574 587 570 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=34260 $D=0
M1575 588 571 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=38890 $D=0
M1576 585 570 580 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=34260 $D=0
M1577 586 571 126 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=38890 $D=0
M1578 581 587 585 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=34260 $D=0
M1579 582 588 586 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=38890 $D=0
M1580 589 583 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=34260 $D=0
M1581 590 584 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=38890 $D=0
M1582 127 583 578 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=34260 $D=0
M1583 580 584 579 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=38890 $D=0
M1584 570 589 127 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=34260 $D=0
M1585 571 590 580 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=38890 $D=0
M1586 591 127 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=34260 $D=0
M1587 592 580 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=38890 $D=0
M1588 593 583 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=34260 $D=0
M1589 594 584 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=38890 $D=0
M1590 595 583 591 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=34260 $D=0
M1591 596 584 592 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=38890 $D=0
M1592 578 593 595 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=34260 $D=0
M1593 579 594 596 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=38890 $D=0
M1594 792 570 9 9 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=33900 $D=0
M1595 793 571 9 9 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=38530 $D=0
M1596 597 578 792 9 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=33900 $D=0
M1597 598 579 793 9 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=38530 $D=0
M1598 599 595 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=34260 $D=0
M1599 600 596 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=38890 $D=0
M1600 601 570 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=34260 $D=0
M1601 602 571 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=38890 $D=0
M1602 9 578 601 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=34260 $D=0
M1603 9 579 602 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=38890 $D=0
M1604 603 570 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=34260 $D=0
M1605 604 571 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=38890 $D=0
M1606 9 578 603 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=34260 $D=0
M1607 9 579 604 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=38890 $D=0
M1608 794 570 9 9 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=34080 $D=0
M1609 795 571 9 9 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=38710 $D=0
M1610 607 578 794 9 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=34080 $D=0
M1611 608 579 795 9 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=38710 $D=0
M1612 9 603 607 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=34260 $D=0
M1613 9 604 608 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=38890 $D=0
M1614 609 130 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=34260 $D=0
M1615 610 130 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=38890 $D=0
M1616 611 130 597 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=34260 $D=0
M1617 612 130 598 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=38890 $D=0
M1618 601 609 611 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=34260 $D=0
M1619 602 610 612 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=38890 $D=0
M1620 613 130 599 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=34260 $D=0
M1621 614 130 600 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=38890 $D=0
M1622 607 609 613 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=34260 $D=0
M1623 608 610 614 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=38890 $D=0
M1624 615 131 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=34260 $D=0
M1625 616 131 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=38890 $D=0
M1626 617 131 613 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=34260 $D=0
M1627 618 131 614 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=38890 $D=0
M1628 611 615 617 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=34260 $D=0
M1629 612 616 618 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=38890 $D=0
M1630 13 617 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=34260 $D=0
M1631 14 618 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=38890 $D=0
M1632 619 132 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=34260 $D=0
M1633 620 132 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=38890 $D=0
M1634 621 132 133 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=34260 $D=0
M1635 622 132 134 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=38890 $D=0
M1636 135 619 621 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=34260 $D=0
M1637 136 620 622 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=38890 $D=0
M1638 623 132 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=34260 $D=0
M1639 624 132 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=38890 $D=0
M1640 625 132 137 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=34260 $D=0
M1641 626 132 138 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=38890 $D=0
M1642 139 623 625 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=34260 $D=0
M1643 140 624 626 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=38890 $D=0
M1644 627 132 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=34260 $D=0
M1645 628 132 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=38890 $D=0
M1646 629 132 128 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=34260 $D=0
M1647 630 132 129 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=38890 $D=0
M1648 141 627 629 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=34260 $D=0
M1649 108 628 630 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=38890 $D=0
M1650 631 132 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=34260 $D=0
M1651 632 132 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=38890 $D=0
M1652 633 132 142 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=34260 $D=0
M1653 634 132 143 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=38890 $D=0
M1654 144 631 633 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=34260 $D=0
M1655 145 632 634 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=38890 $D=0
M1656 635 132 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=34260 $D=0
M1657 636 132 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=38890 $D=0
M1658 637 132 146 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=34260 $D=0
M1659 638 132 147 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=38890 $D=0
M1660 144 635 637 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=34260 $D=0
M1661 144 636 638 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=38890 $D=0
M1662 9 570 782 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=34260 $D=0
M1663 9 571 783 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=38890 $D=0
M1664 136 782 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=34260 $D=0
M1665 133 783 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=38890 $D=0
M1666 639 148 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=34260 $D=0
M1667 640 148 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=38890 $D=0
M1668 149 148 136 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=34260 $D=0
M1669 150 148 133 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=38890 $D=0
M1670 621 639 149 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=34260 $D=0
M1671 622 640 150 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=38890 $D=0
M1672 641 151 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=34260 $D=0
M1673 642 151 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=38890 $D=0
M1674 152 151 149 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=34260 $D=0
M1675 113 151 150 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=38890 $D=0
M1676 625 641 152 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=34260 $D=0
M1677 626 642 113 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=38890 $D=0
M1678 643 153 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=34260 $D=0
M1679 644 153 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=38890 $D=0
M1680 154 153 152 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=34260 $D=0
M1681 106 153 113 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=38890 $D=0
M1682 629 643 154 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=34260 $D=0
M1683 630 644 106 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=38890 $D=0
M1684 645 155 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=34260 $D=0
M1685 646 155 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=38890 $D=0
M1686 156 155 154 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=34260 $D=0
M1687 157 155 106 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=38890 $D=0
M1688 633 645 156 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=34260 $D=0
M1689 634 646 157 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=38890 $D=0
M1690 647 158 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=34260 $D=0
M1691 648 158 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=38890 $D=0
M1692 220 158 156 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=34260 $D=0
M1693 221 158 157 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=38890 $D=0
M1694 637 647 220 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=34260 $D=0
M1695 638 648 221 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=38890 $D=0
M1696 649 159 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=34260 $D=0
M1697 650 159 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=38890 $D=0
M1698 651 159 119 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=34260 $D=0
M1699 652 159 120 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=38890 $D=0
M1700 11 649 651 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=34260 $D=0
M1701 12 650 652 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=38890 $D=0
M1702 653 560 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=34260 $D=0
M1703 654 561 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=38890 $D=0
M1704 9 651 653 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=34260 $D=0
M1705 9 652 654 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=38890 $D=0
M1706 796 560 9 9 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=34080 $D=0
M1707 797 561 9 9 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=38710 $D=0
M1708 657 651 796 9 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=34080 $D=0
M1709 658 652 797 9 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=38710 $D=0
M1710 9 653 657 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=34260 $D=0
M1711 9 654 658 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=38890 $D=0
M1712 784 160 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=34260 $D=0
M1713 785 659 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=38890 $D=0
M1714 9 657 784 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=34260 $D=0
M1715 9 658 785 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=38890 $D=0
M1716 659 784 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=34260 $D=0
M1717 161 785 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=38890 $D=0
M1718 798 560 9 9 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=33900 $D=0
M1719 799 561 9 9 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=38530 $D=0
M1720 660 662 798 9 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=33900 $D=0
M1721 661 663 799 9 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=38530 $D=0
M1722 662 651 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=34260 $D=0
M1723 663 652 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=38890 $D=0
M1724 664 660 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=34260 $D=0
M1725 665 661 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=38890 $D=0
M1726 9 160 664 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=34260 $D=0
M1727 9 659 665 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=38890 $D=0
M1728 667 162 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=34260 $D=0
M1729 668 666 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=38890 $D=0
M1730 666 664 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=34260 $D=0
M1731 163 665 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=38890 $D=0
M1732 9 667 666 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=34260 $D=0
M1733 9 668 163 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=38890 $D=0
M1734 670 669 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=34260 $D=0
M1735 671 164 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=38890 $D=0
M1736 9 674 672 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=34260 $D=0
M1737 9 675 673 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=38890 $D=0
M1738 676 122 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=34260 $D=0
M1739 677 123 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=38890 $D=0
M1740 674 122 669 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=34260 $D=0
M1741 675 123 164 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=38890 $D=0
M1742 670 676 674 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=34260 $D=0
M1743 671 677 675 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=38890 $D=0
M1744 678 672 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=34260 $D=0
M1745 679 673 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=38890 $D=0
M1746 165 672 6 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=34260 $D=0
M1747 669 673 6 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=38890 $D=0
M1748 122 678 165 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=34260 $D=0
M1749 123 679 669 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=38890 $D=0
M1750 680 165 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=34260 $D=0
M1751 681 669 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=38890 $D=0
M1752 682 672 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=34260 $D=0
M1753 683 673 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=38890 $D=0
M1754 222 672 680 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=34260 $D=0
M1755 223 673 681 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=38890 $D=0
M1756 6 682 222 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=34260 $D=0
M1757 6 683 223 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=38890 $D=0
M1758 684 166 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=34260 $D=0
M1759 685 166 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=38890 $D=0
M1760 686 166 222 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=34260 $D=0
M1761 687 166 223 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=38890 $D=0
M1762 13 684 686 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=34260 $D=0
M1763 14 685 687 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=38890 $D=0
M1764 688 167 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=34260 $D=0
M1765 689 167 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=38890 $D=0
M1766 690 167 686 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=34260 $D=0
M1767 691 167 687 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=38890 $D=0
M1768 6 688 690 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=34260 $D=0
M1769 6 689 691 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=38890 $D=0
M1770 692 118 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=34260 $D=0
M1771 693 118 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=38890 $D=0
M1772 9 692 694 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=34260 $D=0
M1773 9 693 695 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=38890 $D=0
M1774 696 118 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=34260 $D=0
M1775 697 118 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=38890 $D=0
M1776 698 694 690 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=34260 $D=0
M1777 699 695 691 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=38890 $D=0
M1778 9 698 786 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=34260 $D=0
M1779 9 699 787 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=38890 $D=0
M1780 700 786 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=34260 $D=0
M1781 701 787 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=38890 $D=0
M1782 698 692 700 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=34260 $D=0
M1783 699 693 701 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=38890 $D=0
M1784 702 696 700 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=34260 $D=0
M1785 703 697 701 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=38890 $D=0
M1786 9 706 704 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=34260 $D=0
M1787 9 707 705 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=38890 $D=0
M1788 706 118 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=34260 $D=0
M1789 707 118 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=38890 $D=0
M1790 788 702 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=34260 $D=0
M1791 789 703 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=38890 $D=0
M1792 708 706 788 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=34260 $D=0
M1793 709 707 789 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=38890 $D=0
M1794 9 708 122 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=34260 $D=0
M1795 9 709 123 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=38890 $D=0
M1796 790 122 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=34260 $D=0
M1797 791 123 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=38890 $D=0
M1798 708 704 790 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=34260 $D=0
M1799 709 705 791 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=38890 $D=0
.ENDS
***************************************
.SUBCKT ICV_39 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 111 112 113 114 115 117 118 119 120 121 122
+ 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 142 143
+ 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162 163
+ 164 165 166
** N=805 EP=163 IP=1514 FDC=1800
M0 190 1 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=23750 $D=1
M1 191 1 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=28380 $D=1
M2 192 190 2 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=23750 $D=1
M3 193 191 3 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=28380 $D=1
M4 6 1 192 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=23750 $D=1
M5 6 1 193 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=28380 $D=1
M6 194 190 4 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=23750 $D=1
M7 195 191 4 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=28380 $D=1
M8 5 1 194 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=23750 $D=1
M9 5 1 195 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=28380 $D=1
M10 196 190 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=23750 $D=1
M11 197 191 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=28380 $D=1
M12 6 1 196 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=23750 $D=1
M13 6 1 197 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=28380 $D=1
M14 200 198 196 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=23750 $D=1
M15 201 199 197 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=28380 $D=1
M16 198 7 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=23750 $D=1
M17 199 7 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=28380 $D=1
M18 202 198 194 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=23750 $D=1
M19 203 199 195 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=28380 $D=1
M20 192 7 202 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=23750 $D=1
M21 193 7 203 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=28380 $D=1
M22 204 8 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=23750 $D=1
M23 205 8 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=28380 $D=1
M24 206 204 202 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=23750 $D=1
M25 207 205 203 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=28380 $D=1
M26 200 8 206 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=23750 $D=1
M27 201 8 207 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=28380 $D=1
M28 208 10 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=23750 $D=1
M29 209 10 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=28380 $D=1
M30 210 208 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=23750 $D=1
M31 211 209 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=28380 $D=1
M32 11 10 210 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=23750 $D=1
M33 12 10 211 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=28380 $D=1
M34 212 208 13 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=23750 $D=1
M35 213 209 14 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=28380 $D=1
M36 214 10 212 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=23750 $D=1
M37 215 10 213 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=28380 $D=1
M38 218 208 216 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=23750 $D=1
M39 219 209 217 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=28380 $D=1
M40 206 10 218 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=23750 $D=1
M41 207 10 219 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=28380 $D=1
M42 222 220 218 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=23750 $D=1
M43 223 221 219 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=28380 $D=1
M44 220 15 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=23750 $D=1
M45 221 15 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=28380 $D=1
M46 224 220 212 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=23750 $D=1
M47 225 221 213 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=28380 $D=1
M48 210 15 224 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=23750 $D=1
M49 211 15 225 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=28380 $D=1
M50 226 16 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=23750 $D=1
M51 227 16 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=28380 $D=1
M52 228 226 224 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=23750 $D=1
M53 229 227 225 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=28380 $D=1
M54 222 16 228 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=23750 $D=1
M55 223 16 229 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=28380 $D=1
M56 6 17 230 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=23750 $D=1
M57 6 17 231 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=28380 $D=1
M58 232 18 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=23750 $D=1
M59 233 18 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=28380 $D=1
M60 234 17 228 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=23750 $D=1
M61 235 17 229 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=28380 $D=1
M62 6 234 704 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=23750 $D=1
M63 6 235 705 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=28380 $D=1
M64 236 704 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=23750 $D=1
M65 237 705 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=28380 $D=1
M66 234 230 236 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=23750 $D=1
M67 235 231 237 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=28380 $D=1
M68 236 18 238 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=23750 $D=1
M69 237 18 239 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=28380 $D=1
M70 242 19 236 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=23750 $D=1
M71 243 19 237 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=28380 $D=1
M72 240 19 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=23750 $D=1
M73 241 19 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=28380 $D=1
M74 6 20 244 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=23750 $D=1
M75 6 20 245 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=28380 $D=1
M76 246 21 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=23750 $D=1
M77 247 21 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=28380 $D=1
M78 248 20 228 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=23750 $D=1
M79 249 20 229 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=28380 $D=1
M80 6 248 706 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=23750 $D=1
M81 6 249 707 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=28380 $D=1
M82 250 706 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=23750 $D=1
M83 251 707 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=28380 $D=1
M84 248 244 250 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=23750 $D=1
M85 249 245 251 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=28380 $D=1
M86 250 21 238 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=23750 $D=1
M87 251 21 239 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=28380 $D=1
M88 242 22 250 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=23750 $D=1
M89 243 22 251 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=28380 $D=1
M90 252 22 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=23750 $D=1
M91 253 22 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=28380 $D=1
M92 6 23 254 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=23750 $D=1
M93 6 23 255 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=28380 $D=1
M94 256 24 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=23750 $D=1
M95 257 24 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=28380 $D=1
M96 258 23 228 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=23750 $D=1
M97 259 23 229 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=28380 $D=1
M98 6 258 708 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=23750 $D=1
M99 6 259 709 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=28380 $D=1
M100 260 708 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=23750 $D=1
M101 261 709 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=28380 $D=1
M102 258 254 260 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=23750 $D=1
M103 259 255 261 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=28380 $D=1
M104 260 24 238 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=23750 $D=1
M105 261 24 239 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=28380 $D=1
M106 242 25 260 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=23750 $D=1
M107 243 25 261 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=28380 $D=1
M108 262 25 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=23750 $D=1
M109 263 25 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=28380 $D=1
M110 6 26 264 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=23750 $D=1
M111 6 26 265 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=28380 $D=1
M112 266 27 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=23750 $D=1
M113 267 27 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=28380 $D=1
M114 268 26 228 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=23750 $D=1
M115 269 26 229 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=28380 $D=1
M116 6 268 710 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=23750 $D=1
M117 6 269 711 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=28380 $D=1
M118 270 710 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=23750 $D=1
M119 271 711 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=28380 $D=1
M120 268 264 270 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=23750 $D=1
M121 269 265 271 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=28380 $D=1
M122 270 27 238 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=23750 $D=1
M123 271 27 239 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=28380 $D=1
M124 242 28 270 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=23750 $D=1
M125 243 28 271 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=28380 $D=1
M126 272 28 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=23750 $D=1
M127 273 28 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=28380 $D=1
M128 6 29 274 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=23750 $D=1
M129 6 29 275 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=28380 $D=1
M130 276 30 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=23750 $D=1
M131 277 30 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=28380 $D=1
M132 278 29 228 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=23750 $D=1
M133 279 29 229 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=28380 $D=1
M134 6 278 712 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=23750 $D=1
M135 6 279 713 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=28380 $D=1
M136 280 712 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=23750 $D=1
M137 281 713 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=28380 $D=1
M138 278 274 280 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=23750 $D=1
M139 279 275 281 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=28380 $D=1
M140 280 30 238 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=23750 $D=1
M141 281 30 239 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=28380 $D=1
M142 242 31 280 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=23750 $D=1
M143 243 31 281 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=28380 $D=1
M144 282 31 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=23750 $D=1
M145 283 31 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=28380 $D=1
M146 6 32 284 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=23750 $D=1
M147 6 32 285 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=28380 $D=1
M148 286 33 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=23750 $D=1
M149 287 33 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=28380 $D=1
M150 288 32 228 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=23750 $D=1
M151 289 32 229 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=28380 $D=1
M152 6 288 714 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=23750 $D=1
M153 6 289 715 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=28380 $D=1
M154 290 714 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=23750 $D=1
M155 291 715 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=28380 $D=1
M156 288 284 290 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=23750 $D=1
M157 289 285 291 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=28380 $D=1
M158 290 33 238 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=23750 $D=1
M159 291 33 239 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=28380 $D=1
M160 242 34 290 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=23750 $D=1
M161 243 34 291 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=28380 $D=1
M162 292 34 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=23750 $D=1
M163 293 34 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=28380 $D=1
M164 6 35 294 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=23750 $D=1
M165 6 35 295 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=28380 $D=1
M166 296 36 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=23750 $D=1
M167 297 36 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=28380 $D=1
M168 298 35 228 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=23750 $D=1
M169 299 35 229 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=28380 $D=1
M170 6 298 716 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=23750 $D=1
M171 6 299 717 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=28380 $D=1
M172 300 716 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=23750 $D=1
M173 301 717 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=28380 $D=1
M174 298 294 300 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=23750 $D=1
M175 299 295 301 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=28380 $D=1
M176 300 36 238 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=23750 $D=1
M177 301 36 239 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=28380 $D=1
M178 242 37 300 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=23750 $D=1
M179 243 37 301 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=28380 $D=1
M180 302 37 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=23750 $D=1
M181 303 37 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=28380 $D=1
M182 6 38 304 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=23750 $D=1
M183 6 38 305 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=28380 $D=1
M184 306 39 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=23750 $D=1
M185 307 39 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=28380 $D=1
M186 308 38 228 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=23750 $D=1
M187 309 38 229 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=28380 $D=1
M188 6 308 718 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=23750 $D=1
M189 6 309 719 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=28380 $D=1
M190 310 718 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=23750 $D=1
M191 311 719 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=28380 $D=1
M192 308 304 310 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=23750 $D=1
M193 309 305 311 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=28380 $D=1
M194 310 39 238 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=23750 $D=1
M195 311 39 239 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=28380 $D=1
M196 242 40 310 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=23750 $D=1
M197 243 40 311 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=28380 $D=1
M198 312 40 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=23750 $D=1
M199 313 40 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=28380 $D=1
M200 6 41 314 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=23750 $D=1
M201 6 41 315 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=28380 $D=1
M202 316 42 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=23750 $D=1
M203 317 42 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=28380 $D=1
M204 318 41 228 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=23750 $D=1
M205 319 41 229 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=28380 $D=1
M206 6 318 720 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=23750 $D=1
M207 6 319 721 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=28380 $D=1
M208 320 720 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=23750 $D=1
M209 321 721 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=28380 $D=1
M210 318 314 320 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=23750 $D=1
M211 319 315 321 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=28380 $D=1
M212 320 42 238 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=23750 $D=1
M213 321 42 239 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=28380 $D=1
M214 242 43 320 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=23750 $D=1
M215 243 43 321 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=28380 $D=1
M216 322 43 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=23750 $D=1
M217 323 43 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=28380 $D=1
M218 6 44 324 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=23750 $D=1
M219 6 44 325 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=28380 $D=1
M220 326 45 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=23750 $D=1
M221 327 45 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=28380 $D=1
M222 328 44 228 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=23750 $D=1
M223 329 44 229 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=28380 $D=1
M224 6 328 722 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=23750 $D=1
M225 6 329 723 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=28380 $D=1
M226 330 722 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=23750 $D=1
M227 331 723 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=28380 $D=1
M228 328 324 330 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=23750 $D=1
M229 329 325 331 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=28380 $D=1
M230 330 45 238 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=23750 $D=1
M231 331 45 239 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=28380 $D=1
M232 242 46 330 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=23750 $D=1
M233 243 46 331 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=28380 $D=1
M234 332 46 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=23750 $D=1
M235 333 46 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=28380 $D=1
M236 6 47 334 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=23750 $D=1
M237 6 47 335 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=28380 $D=1
M238 336 48 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=23750 $D=1
M239 337 48 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=28380 $D=1
M240 338 47 228 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=23750 $D=1
M241 339 47 229 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=28380 $D=1
M242 6 338 724 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=23750 $D=1
M243 6 339 725 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=28380 $D=1
M244 340 724 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=23750 $D=1
M245 341 725 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=28380 $D=1
M246 338 334 340 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=23750 $D=1
M247 339 335 341 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=28380 $D=1
M248 340 48 238 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=23750 $D=1
M249 341 48 239 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=28380 $D=1
M250 242 49 340 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=23750 $D=1
M251 243 49 341 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=28380 $D=1
M252 342 49 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=23750 $D=1
M253 343 49 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=28380 $D=1
M254 6 50 344 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=23750 $D=1
M255 6 50 345 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=28380 $D=1
M256 346 51 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=23750 $D=1
M257 347 51 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=28380 $D=1
M258 348 50 228 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=23750 $D=1
M259 349 50 229 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=28380 $D=1
M260 6 348 726 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=23750 $D=1
M261 6 349 727 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=28380 $D=1
M262 350 726 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=23750 $D=1
M263 351 727 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=28380 $D=1
M264 348 344 350 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=23750 $D=1
M265 349 345 351 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=28380 $D=1
M266 350 51 238 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=23750 $D=1
M267 351 51 239 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=28380 $D=1
M268 242 52 350 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=23750 $D=1
M269 243 52 351 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=28380 $D=1
M270 352 52 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=23750 $D=1
M271 353 52 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=28380 $D=1
M272 6 53 354 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=23750 $D=1
M273 6 53 355 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=28380 $D=1
M274 356 54 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=23750 $D=1
M275 357 54 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=28380 $D=1
M276 358 53 228 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=23750 $D=1
M277 359 53 229 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=28380 $D=1
M278 6 358 728 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=23750 $D=1
M279 6 359 729 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=28380 $D=1
M280 360 728 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=23750 $D=1
M281 361 729 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=28380 $D=1
M282 358 354 360 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=23750 $D=1
M283 359 355 361 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=28380 $D=1
M284 360 54 238 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=23750 $D=1
M285 361 54 239 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=28380 $D=1
M286 242 55 360 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=23750 $D=1
M287 243 55 361 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=28380 $D=1
M288 362 55 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=23750 $D=1
M289 363 55 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=28380 $D=1
M290 6 56 364 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=23750 $D=1
M291 6 56 365 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=28380 $D=1
M292 366 57 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=23750 $D=1
M293 367 57 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=28380 $D=1
M294 368 56 228 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=23750 $D=1
M295 369 56 229 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=28380 $D=1
M296 6 368 730 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=23750 $D=1
M297 6 369 731 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=28380 $D=1
M298 370 730 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=23750 $D=1
M299 371 731 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=28380 $D=1
M300 368 364 370 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=23750 $D=1
M301 369 365 371 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=28380 $D=1
M302 370 57 238 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=23750 $D=1
M303 371 57 239 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=28380 $D=1
M304 242 58 370 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=23750 $D=1
M305 243 58 371 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=28380 $D=1
M306 372 58 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=23750 $D=1
M307 373 58 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=28380 $D=1
M308 6 59 374 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=23750 $D=1
M309 6 59 375 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=28380 $D=1
M310 376 60 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=23750 $D=1
M311 377 60 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=28380 $D=1
M312 378 59 228 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=23750 $D=1
M313 379 59 229 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=28380 $D=1
M314 6 378 732 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=23750 $D=1
M315 6 379 733 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=28380 $D=1
M316 380 732 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=23750 $D=1
M317 381 733 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=28380 $D=1
M318 378 374 380 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=23750 $D=1
M319 379 375 381 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=28380 $D=1
M320 380 60 238 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=23750 $D=1
M321 381 60 239 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=28380 $D=1
M322 242 61 380 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=23750 $D=1
M323 243 61 381 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=28380 $D=1
M324 382 61 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=23750 $D=1
M325 383 61 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=28380 $D=1
M326 6 62 384 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=23750 $D=1
M327 6 62 385 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=28380 $D=1
M328 386 63 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=23750 $D=1
M329 387 63 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=28380 $D=1
M330 388 62 228 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=23750 $D=1
M331 389 62 229 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=28380 $D=1
M332 6 388 734 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=23750 $D=1
M333 6 389 735 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=28380 $D=1
M334 390 734 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=23750 $D=1
M335 391 735 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=28380 $D=1
M336 388 384 390 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=23750 $D=1
M337 389 385 391 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=28380 $D=1
M338 390 63 238 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=23750 $D=1
M339 391 63 239 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=28380 $D=1
M340 242 64 390 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=23750 $D=1
M341 243 64 391 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=28380 $D=1
M342 392 64 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=23750 $D=1
M343 393 64 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=28380 $D=1
M344 6 65 394 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=23750 $D=1
M345 6 65 395 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=28380 $D=1
M346 396 66 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=23750 $D=1
M347 397 66 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=28380 $D=1
M348 398 65 228 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=23750 $D=1
M349 399 65 229 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=28380 $D=1
M350 6 398 736 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=23750 $D=1
M351 6 399 737 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=28380 $D=1
M352 400 736 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=23750 $D=1
M353 401 737 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=28380 $D=1
M354 398 394 400 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=23750 $D=1
M355 399 395 401 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=28380 $D=1
M356 400 66 238 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=23750 $D=1
M357 401 66 239 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=28380 $D=1
M358 242 67 400 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=23750 $D=1
M359 243 67 401 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=28380 $D=1
M360 402 67 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=23750 $D=1
M361 403 67 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=28380 $D=1
M362 6 68 404 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=23750 $D=1
M363 6 68 405 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=28380 $D=1
M364 406 69 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=23750 $D=1
M365 407 69 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=28380 $D=1
M366 408 68 228 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=23750 $D=1
M367 409 68 229 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=28380 $D=1
M368 6 408 738 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=23750 $D=1
M369 6 409 739 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=28380 $D=1
M370 410 738 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=23750 $D=1
M371 411 739 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=28380 $D=1
M372 408 404 410 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=23750 $D=1
M373 409 405 411 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=28380 $D=1
M374 410 69 238 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=23750 $D=1
M375 411 69 239 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=28380 $D=1
M376 242 70 410 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=23750 $D=1
M377 243 70 411 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=28380 $D=1
M378 412 70 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=23750 $D=1
M379 413 70 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=28380 $D=1
M380 6 71 414 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=23750 $D=1
M381 6 71 415 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=28380 $D=1
M382 416 72 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=23750 $D=1
M383 417 72 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=28380 $D=1
M384 418 71 228 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=23750 $D=1
M385 419 71 229 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=28380 $D=1
M386 6 418 740 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=23750 $D=1
M387 6 419 741 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=28380 $D=1
M388 420 740 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=23750 $D=1
M389 421 741 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=28380 $D=1
M390 418 414 420 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=23750 $D=1
M391 419 415 421 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=28380 $D=1
M392 420 72 238 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=23750 $D=1
M393 421 72 239 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=28380 $D=1
M394 242 73 420 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=23750 $D=1
M395 243 73 421 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=28380 $D=1
M396 422 73 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=23750 $D=1
M397 423 73 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=28380 $D=1
M398 6 74 424 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=23750 $D=1
M399 6 74 425 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=28380 $D=1
M400 426 75 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=23750 $D=1
M401 427 75 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=28380 $D=1
M402 428 74 228 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=23750 $D=1
M403 429 74 229 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=28380 $D=1
M404 6 428 742 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=23750 $D=1
M405 6 429 743 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=28380 $D=1
M406 430 742 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=23750 $D=1
M407 431 743 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=28380 $D=1
M408 428 424 430 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=23750 $D=1
M409 429 425 431 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=28380 $D=1
M410 430 75 238 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=23750 $D=1
M411 431 75 239 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=28380 $D=1
M412 242 76 430 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=23750 $D=1
M413 243 76 431 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=28380 $D=1
M414 432 76 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=23750 $D=1
M415 433 76 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=28380 $D=1
M416 6 77 434 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=23750 $D=1
M417 6 77 435 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=28380 $D=1
M418 436 78 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=23750 $D=1
M419 437 78 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=28380 $D=1
M420 438 77 228 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=23750 $D=1
M421 439 77 229 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=28380 $D=1
M422 6 438 744 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=23750 $D=1
M423 6 439 745 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=28380 $D=1
M424 440 744 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=23750 $D=1
M425 441 745 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=28380 $D=1
M426 438 434 440 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=23750 $D=1
M427 439 435 441 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=28380 $D=1
M428 440 78 238 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=23750 $D=1
M429 441 78 239 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=28380 $D=1
M430 242 79 440 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=23750 $D=1
M431 243 79 441 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=28380 $D=1
M432 442 79 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=23750 $D=1
M433 443 79 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=28380 $D=1
M434 6 80 444 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=23750 $D=1
M435 6 80 445 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=28380 $D=1
M436 446 81 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=23750 $D=1
M437 447 81 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=28380 $D=1
M438 448 80 228 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=23750 $D=1
M439 449 80 229 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=28380 $D=1
M440 6 448 746 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=23750 $D=1
M441 6 449 747 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=28380 $D=1
M442 450 746 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=23750 $D=1
M443 451 747 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=28380 $D=1
M444 448 444 450 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=23750 $D=1
M445 449 445 451 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=28380 $D=1
M446 450 81 238 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=23750 $D=1
M447 451 81 239 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=28380 $D=1
M448 242 82 450 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=23750 $D=1
M449 243 82 451 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=28380 $D=1
M450 452 82 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=23750 $D=1
M451 453 82 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=28380 $D=1
M452 6 83 454 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=23750 $D=1
M453 6 83 455 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=28380 $D=1
M454 456 84 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=23750 $D=1
M455 457 84 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=28380 $D=1
M456 458 83 228 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=23750 $D=1
M457 459 83 229 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=28380 $D=1
M458 6 458 748 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=23750 $D=1
M459 6 459 749 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=28380 $D=1
M460 460 748 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=23750 $D=1
M461 461 749 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=28380 $D=1
M462 458 454 460 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=23750 $D=1
M463 459 455 461 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=28380 $D=1
M464 460 84 238 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=23750 $D=1
M465 461 84 239 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=28380 $D=1
M466 242 85 460 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=23750 $D=1
M467 243 85 461 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=28380 $D=1
M468 462 85 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=23750 $D=1
M469 463 85 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=28380 $D=1
M470 6 86 464 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=23750 $D=1
M471 6 86 465 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=28380 $D=1
M472 466 87 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=23750 $D=1
M473 467 87 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=28380 $D=1
M474 468 86 228 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=23750 $D=1
M475 469 86 229 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=28380 $D=1
M476 6 468 750 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=23750 $D=1
M477 6 469 751 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=28380 $D=1
M478 470 750 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=23750 $D=1
M479 471 751 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=28380 $D=1
M480 468 464 470 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=23750 $D=1
M481 469 465 471 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=28380 $D=1
M482 470 87 238 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=23750 $D=1
M483 471 87 239 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=28380 $D=1
M484 242 88 470 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=23750 $D=1
M485 243 88 471 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=28380 $D=1
M486 472 88 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=23750 $D=1
M487 473 88 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=28380 $D=1
M488 6 89 474 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=23750 $D=1
M489 6 89 475 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=28380 $D=1
M490 476 90 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=23750 $D=1
M491 477 90 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=28380 $D=1
M492 478 89 228 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=23750 $D=1
M493 479 89 229 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=28380 $D=1
M494 6 478 752 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=23750 $D=1
M495 6 479 753 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=28380 $D=1
M496 480 752 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=23750 $D=1
M497 481 753 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=28380 $D=1
M498 478 474 480 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=23750 $D=1
M499 479 475 481 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=28380 $D=1
M500 480 90 238 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=23750 $D=1
M501 481 90 239 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=28380 $D=1
M502 242 91 480 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=23750 $D=1
M503 243 91 481 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=28380 $D=1
M504 482 91 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=23750 $D=1
M505 483 91 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=28380 $D=1
M506 6 92 484 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=23750 $D=1
M507 6 92 485 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=28380 $D=1
M508 486 93 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=23750 $D=1
M509 487 93 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=28380 $D=1
M510 488 92 228 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=23750 $D=1
M511 489 92 229 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=28380 $D=1
M512 6 488 754 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=23750 $D=1
M513 6 489 755 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=28380 $D=1
M514 490 754 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=23750 $D=1
M515 491 755 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=28380 $D=1
M516 488 484 490 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=23750 $D=1
M517 489 485 491 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=28380 $D=1
M518 490 93 238 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=23750 $D=1
M519 491 93 239 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=28380 $D=1
M520 242 94 490 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=23750 $D=1
M521 243 94 491 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=28380 $D=1
M522 492 94 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=23750 $D=1
M523 493 94 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=28380 $D=1
M524 6 95 494 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=23750 $D=1
M525 6 95 495 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=28380 $D=1
M526 496 96 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=23750 $D=1
M527 497 96 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=28380 $D=1
M528 498 95 228 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=23750 $D=1
M529 499 95 229 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=28380 $D=1
M530 6 498 756 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=23750 $D=1
M531 6 499 757 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=28380 $D=1
M532 500 756 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=23750 $D=1
M533 501 757 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=28380 $D=1
M534 498 494 500 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=23750 $D=1
M535 499 495 501 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=28380 $D=1
M536 500 96 238 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=23750 $D=1
M537 501 96 239 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=28380 $D=1
M538 242 97 500 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=23750 $D=1
M539 243 97 501 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=28380 $D=1
M540 502 97 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=23750 $D=1
M541 503 97 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=28380 $D=1
M542 6 98 504 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=23750 $D=1
M543 6 98 505 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=28380 $D=1
M544 506 99 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=23750 $D=1
M545 507 99 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=28380 $D=1
M546 508 98 228 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=23750 $D=1
M547 509 98 229 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=28380 $D=1
M548 6 508 758 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=23750 $D=1
M549 6 509 759 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=28380 $D=1
M550 510 758 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=23750 $D=1
M551 511 759 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=28380 $D=1
M552 508 504 510 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=23750 $D=1
M553 509 505 511 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=28380 $D=1
M554 510 99 238 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=23750 $D=1
M555 511 99 239 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=28380 $D=1
M556 242 100 510 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=23750 $D=1
M557 243 100 511 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=28380 $D=1
M558 512 100 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=23750 $D=1
M559 513 100 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=28380 $D=1
M560 6 101 514 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=23750 $D=1
M561 6 101 515 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=28380 $D=1
M562 516 102 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=23750 $D=1
M563 517 102 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=28380 $D=1
M564 518 101 228 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=23750 $D=1
M565 519 101 229 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=28380 $D=1
M566 6 518 760 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=23750 $D=1
M567 6 519 761 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=28380 $D=1
M568 520 760 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=23750 $D=1
M569 521 761 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=28380 $D=1
M570 518 514 520 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=23750 $D=1
M571 519 515 521 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=28380 $D=1
M572 520 102 238 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=23750 $D=1
M573 521 102 239 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=28380 $D=1
M574 242 103 520 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=23750 $D=1
M575 243 103 521 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=28380 $D=1
M576 522 103 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=23750 $D=1
M577 523 103 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=28380 $D=1
M578 6 104 524 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=23750 $D=1
M579 6 104 525 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=28380 $D=1
M580 526 105 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=23750 $D=1
M581 527 105 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=28380 $D=1
M582 528 104 228 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=23750 $D=1
M583 529 104 229 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=28380 $D=1
M584 6 528 762 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=23750 $D=1
M585 6 529 763 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=28380 $D=1
M586 530 762 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=23750 $D=1
M587 531 763 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=28380 $D=1
M588 528 524 530 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=23750 $D=1
M589 529 525 531 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=28380 $D=1
M590 530 105 238 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=23750 $D=1
M591 531 105 239 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=28380 $D=1
M592 242 107 530 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=23750 $D=1
M593 243 107 531 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=28380 $D=1
M594 532 107 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=23750 $D=1
M595 533 107 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=28380 $D=1
M596 6 108 534 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=23750 $D=1
M597 6 108 535 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=28380 $D=1
M598 536 109 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=23750 $D=1
M599 537 109 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=28380 $D=1
M600 538 108 228 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=23750 $D=1
M601 539 108 229 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=28380 $D=1
M602 6 538 764 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=23750 $D=1
M603 6 539 765 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=28380 $D=1
M604 540 764 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=23750 $D=1
M605 541 765 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=28380 $D=1
M606 538 534 540 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=23750 $D=1
M607 539 535 541 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=28380 $D=1
M608 540 109 238 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=23750 $D=1
M609 541 109 239 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=28380 $D=1
M610 242 111 540 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=23750 $D=1
M611 243 111 541 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=28380 $D=1
M612 542 111 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=23750 $D=1
M613 543 111 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=28380 $D=1
M614 6 112 544 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=23750 $D=1
M615 6 112 545 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=28380 $D=1
M616 546 113 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=23750 $D=1
M617 547 113 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=28380 $D=1
M618 6 113 238 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=23750 $D=1
M619 6 113 239 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=28380 $D=1
M620 242 112 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=23750 $D=1
M621 243 112 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=28380 $D=1
M622 6 550 548 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=23750 $D=1
M623 6 551 549 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=28380 $D=1
M624 550 115 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=23750 $D=1
M625 551 115 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=28380 $D=1
M626 766 238 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=23750 $D=1
M627 767 239 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=28380 $D=1
M628 552 548 766 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=23750 $D=1
M629 553 549 767 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=28380 $D=1
M630 6 552 554 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=23750 $D=1
M631 6 553 555 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=28380 $D=1
M632 768 554 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=23750 $D=1
M633 769 555 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=28380 $D=1
M634 552 550 768 6 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=23750 $D=1
M635 553 551 769 6 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=28380 $D=1
M636 6 558 556 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=23750 $D=1
M637 6 559 557 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=28380 $D=1
M638 558 115 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=23750 $D=1
M639 559 115 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=28380 $D=1
M640 770 242 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=23750 $D=1
M641 771 243 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=28380 $D=1
M642 560 556 770 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=23750 $D=1
M643 561 557 771 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=28380 $D=1
M644 6 560 117 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=23750 $D=1
M645 6 561 118 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=28380 $D=1
M646 772 117 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=23750 $D=1
M647 773 118 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=28380 $D=1
M648 560 558 772 6 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=23750 $D=1
M649 561 559 773 6 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=28380 $D=1
M650 562 119 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=23750 $D=1
M651 563 119 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=28380 $D=1
M652 564 562 554 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=23750 $D=1
M653 565 563 555 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=28380 $D=1
M654 120 119 564 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=23750 $D=1
M655 121 119 565 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=28380 $D=1
M656 566 122 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=23750 $D=1
M657 567 122 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=28380 $D=1
M658 568 566 117 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=23750 $D=1
M659 569 567 118 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=28380 $D=1
M660 774 122 568 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=23750 $D=1
M661 775 122 569 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=28380 $D=1
M662 6 117 774 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=23750 $D=1
M663 6 118 775 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=28380 $D=1
M664 570 123 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=23750 $D=1
M665 571 123 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=28380 $D=1
M666 572 570 568 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=23750 $D=1
M667 573 571 569 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=28380 $D=1
M668 11 123 572 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=23750 $D=1
M669 12 123 573 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=28380 $D=1
M670 575 574 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=23750 $D=1
M671 576 124 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=28380 $D=1
M672 6 579 577 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=23750 $D=1
M673 6 580 578 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=28380 $D=1
M674 581 564 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=23750 $D=1
M675 582 565 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=28380 $D=1
M676 579 581 574 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=23750 $D=1
M677 580 582 124 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=28380 $D=1
M678 575 564 579 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=23750 $D=1
M679 576 565 580 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=28380 $D=1
M680 583 577 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=23750 $D=1
M681 584 578 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=28380 $D=1
M682 125 583 572 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=23750 $D=1
M683 574 584 573 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=28380 $D=1
M684 564 577 125 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=23750 $D=1
M685 565 578 574 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=28380 $D=1
M686 585 125 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=23750 $D=1
M687 586 574 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=28380 $D=1
M688 587 577 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=23750 $D=1
M689 588 578 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=28380 $D=1
M690 589 587 585 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=23750 $D=1
M691 590 588 586 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=28380 $D=1
M692 572 577 589 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=23750 $D=1
M693 573 578 590 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=28380 $D=1
M694 591 564 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=23750 $D=1
M695 592 565 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=28380 $D=1
M696 6 572 591 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=23750 $D=1
M697 6 573 592 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=28380 $D=1
M698 593 589 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=23750 $D=1
M699 594 590 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=28380 $D=1
M700 794 564 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=23750 $D=1
M701 795 565 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=28380 $D=1
M702 595 572 794 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=23750 $D=1
M703 596 573 795 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=28380 $D=1
M704 796 564 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=23750 $D=1
M705 797 565 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=28380 $D=1
M706 597 572 796 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=23750 $D=1
M707 598 573 797 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=28380 $D=1
M708 601 564 599 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=23750 $D=1
M709 602 565 600 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=28380 $D=1
M710 599 572 601 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=23750 $D=1
M711 600 573 602 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=28380 $D=1
M712 6 597 599 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=23750 $D=1
M713 6 598 600 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=28380 $D=1
M714 603 128 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=23750 $D=1
M715 604 128 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=28380 $D=1
M716 605 603 591 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=23750 $D=1
M717 606 604 592 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=28380 $D=1
M718 595 128 605 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=23750 $D=1
M719 596 128 606 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=28380 $D=1
M720 607 603 593 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=23750 $D=1
M721 608 604 594 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=28380 $D=1
M722 601 128 607 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=23750 $D=1
M723 602 128 608 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=28380 $D=1
M724 609 129 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=23750 $D=1
M725 610 129 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=28380 $D=1
M726 611 609 607 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=23750 $D=1
M727 612 610 608 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=28380 $D=1
M728 605 129 611 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=23750 $D=1
M729 606 129 612 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=28380 $D=1
M730 13 611 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=23750 $D=1
M731 14 612 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=28380 $D=1
M732 613 130 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=23750 $D=1
M733 614 130 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=28380 $D=1
M734 615 613 131 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=23750 $D=1
M735 616 614 132 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=28380 $D=1
M736 133 130 615 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=23750 $D=1
M737 134 130 616 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=28380 $D=1
M738 617 130 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=23750 $D=1
M739 618 130 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=28380 $D=1
M740 619 617 135 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=23750 $D=1
M741 620 618 136 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=28380 $D=1
M742 137 130 619 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=23750 $D=1
M743 138 130 620 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=28380 $D=1
M744 621 130 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=23750 $D=1
M745 622 130 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=28380 $D=1
M746 623 621 127 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=23750 $D=1
M747 624 622 126 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=28380 $D=1
M748 139 130 623 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=23750 $D=1
M749 140 130 624 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=28380 $D=1
M750 625 130 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=23750 $D=1
M751 626 130 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=28380 $D=1
M752 627 625 142 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=23750 $D=1
M753 628 626 143 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=28380 $D=1
M754 144 130 627 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=23750 $D=1
M755 144 130 628 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=28380 $D=1
M756 629 130 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=23750 $D=1
M757 630 130 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=28380 $D=1
M758 631 629 145 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=23750 $D=1
M759 632 630 146 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=28380 $D=1
M760 144 130 631 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=23750 $D=1
M761 144 130 632 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=28380 $D=1
M762 6 564 776 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=23750 $D=1
M763 6 565 777 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=28380 $D=1
M764 134 776 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=23750 $D=1
M765 131 777 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=28380 $D=1
M766 633 147 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=23750 $D=1
M767 634 147 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=28380 $D=1
M768 148 633 134 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=23750 $D=1
M769 149 634 131 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=28380 $D=1
M770 615 147 148 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=23750 $D=1
M771 616 147 149 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=28380 $D=1
M772 635 150 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=23750 $D=1
M773 636 150 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=28380 $D=1
M774 151 635 148 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=23750 $D=1
M775 106 636 149 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=28380 $D=1
M776 619 150 151 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=23750 $D=1
M777 620 150 106 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=28380 $D=1
M778 637 152 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=23750 $D=1
M779 638 152 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=28380 $D=1
M780 153 637 151 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=23750 $D=1
M781 114 638 106 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=28380 $D=1
M782 623 152 153 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=23750 $D=1
M783 624 152 114 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=28380 $D=1
M784 639 154 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=23750 $D=1
M785 640 154 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=28380 $D=1
M786 155 639 153 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=23750 $D=1
M787 156 640 114 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=28380 $D=1
M788 627 154 155 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=23750 $D=1
M789 628 154 156 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=28380 $D=1
M790 641 157 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=23750 $D=1
M791 642 157 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=28380 $D=1
M792 214 641 155 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=23750 $D=1
M793 215 642 156 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=28380 $D=1
M794 631 157 214 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=23750 $D=1
M795 632 157 215 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=28380 $D=1
M796 643 158 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=23750 $D=1
M797 644 158 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=28380 $D=1
M798 645 643 117 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=23750 $D=1
M799 646 644 118 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=28380 $D=1
M800 11 158 645 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=23750 $D=1
M801 12 158 646 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=28380 $D=1
M802 798 554 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=23750 $D=1
M803 799 555 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=28380 $D=1
M804 647 645 798 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=23750 $D=1
M805 648 646 799 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=28380 $D=1
M806 651 554 649 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=23750 $D=1
M807 652 555 650 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=28380 $D=1
M808 649 645 651 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=23750 $D=1
M809 650 646 652 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=28380 $D=1
M810 6 647 649 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=23750 $D=1
M811 6 648 650 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=28380 $D=1
M812 800 159 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=23750 $D=1
M813 801 653 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=28380 $D=1
M814 778 651 800 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=23750 $D=1
M815 779 652 801 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=28380 $D=1
M816 653 778 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=23750 $D=1
M817 160 779 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=28380 $D=1
M818 654 554 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=23750 $D=1
M819 655 555 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=28380 $D=1
M820 6 656 654 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=23750 $D=1
M821 6 657 655 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=28380 $D=1
M822 656 645 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=23750 $D=1
M823 657 646 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=28380 $D=1
M824 802 654 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=23750 $D=1
M825 803 655 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=28380 $D=1
M826 658 159 802 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=23750 $D=1
M827 659 653 803 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=28380 $D=1
M828 661 161 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=23750 $D=1
M829 662 660 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=28380 $D=1
M830 804 658 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=23750 $D=1
M831 805 659 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=28380 $D=1
M832 660 661 804 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=23750 $D=1
M833 162 662 805 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=28380 $D=1
M834 664 663 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=23750 $D=1
M835 665 163 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=28380 $D=1
M836 6 668 666 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=23750 $D=1
M837 6 669 667 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=28380 $D=1
M838 670 120 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=23750 $D=1
M839 671 121 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=28380 $D=1
M840 668 670 663 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=23750 $D=1
M841 669 671 163 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=28380 $D=1
M842 664 120 668 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=23750 $D=1
M843 665 121 669 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=28380 $D=1
M844 672 666 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=23750 $D=1
M845 673 667 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=28380 $D=1
M846 164 672 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=23750 $D=1
M847 663 673 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=28380 $D=1
M848 120 666 164 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=23750 $D=1
M849 121 667 663 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=28380 $D=1
M850 674 164 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=23750 $D=1
M851 675 663 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=28380 $D=1
M852 676 666 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=23750 $D=1
M853 677 667 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=28380 $D=1
M854 216 676 674 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=23750 $D=1
M855 217 677 675 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=28380 $D=1
M856 6 666 216 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=23750 $D=1
M857 6 667 217 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=28380 $D=1
M858 678 165 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=23750 $D=1
M859 679 165 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=28380 $D=1
M860 680 678 216 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=23750 $D=1
M861 681 679 217 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=28380 $D=1
M862 13 165 680 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=23750 $D=1
M863 14 165 681 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=28380 $D=1
M864 682 166 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=23750 $D=1
M865 683 166 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=28380 $D=1
M866 684 682 680 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=23750 $D=1
M867 685 683 681 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=28380 $D=1
M868 6 166 684 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=23750 $D=1
M869 6 166 685 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=28380 $D=1
M870 686 115 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=23750 $D=1
M871 687 115 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=28380 $D=1
M872 6 686 688 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=23750 $D=1
M873 6 687 689 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=28380 $D=1
M874 690 115 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=23750 $D=1
M875 691 115 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=28380 $D=1
M876 692 686 684 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=23750 $D=1
M877 693 687 685 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=28380 $D=1
M878 6 692 780 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=23750 $D=1
M879 6 693 781 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=28380 $D=1
M880 694 780 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=23750 $D=1
M881 695 781 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=28380 $D=1
M882 692 688 694 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=23750 $D=1
M883 693 689 695 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=28380 $D=1
M884 696 115 694 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=23750 $D=1
M885 697 115 695 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=28380 $D=1
M886 6 700 698 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=23750 $D=1
M887 6 701 699 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=28380 $D=1
M888 700 115 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=23750 $D=1
M889 701 115 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=28380 $D=1
M890 782 696 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=23750 $D=1
M891 783 697 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=28380 $D=1
M892 702 698 782 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=23750 $D=1
M893 703 699 783 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=28380 $D=1
M894 6 702 120 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=23750 $D=1
M895 6 703 121 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=28380 $D=1
M896 784 120 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=23750 $D=1
M897 785 121 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=28380 $D=1
M898 702 700 784 6 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=23750 $D=1
M899 703 701 785 6 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=28380 $D=1
M900 190 1 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=25000 $D=0
M901 191 1 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=29630 $D=0
M902 192 1 2 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=25000 $D=0
M903 193 1 3 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=29630 $D=0
M904 6 190 192 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=25000 $D=0
M905 6 191 193 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=29630 $D=0
M906 194 1 4 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=25000 $D=0
M907 195 1 4 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=29630 $D=0
M908 5 190 194 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=25000 $D=0
M909 5 191 195 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=29630 $D=0
M910 196 1 6 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=25000 $D=0
M911 197 1 6 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=29630 $D=0
M912 6 190 196 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=25000 $D=0
M913 6 191 197 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=29630 $D=0
M914 200 7 196 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=25000 $D=0
M915 201 7 197 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=29630 $D=0
M916 198 7 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=25000 $D=0
M917 199 7 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=29630 $D=0
M918 202 7 194 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=25000 $D=0
M919 203 7 195 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=29630 $D=0
M920 192 198 202 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=25000 $D=0
M921 193 199 203 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=29630 $D=0
M922 204 8 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=25000 $D=0
M923 205 8 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=29630 $D=0
M924 206 8 202 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=25000 $D=0
M925 207 8 203 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=29630 $D=0
M926 200 204 206 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=25000 $D=0
M927 201 205 207 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=29630 $D=0
M928 208 10 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=25000 $D=0
M929 209 10 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=29630 $D=0
M930 210 10 6 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=25000 $D=0
M931 211 10 6 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=29630 $D=0
M932 11 208 210 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=25000 $D=0
M933 12 209 211 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=29630 $D=0
M934 212 10 13 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=25000 $D=0
M935 213 10 14 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=29630 $D=0
M936 214 208 212 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=25000 $D=0
M937 215 209 213 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=29630 $D=0
M938 218 10 216 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=25000 $D=0
M939 219 10 217 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=29630 $D=0
M940 206 208 218 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=25000 $D=0
M941 207 209 219 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=29630 $D=0
M942 222 15 218 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=25000 $D=0
M943 223 15 219 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=29630 $D=0
M944 220 15 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=25000 $D=0
M945 221 15 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=29630 $D=0
M946 224 15 212 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=25000 $D=0
M947 225 15 213 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=29630 $D=0
M948 210 220 224 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=25000 $D=0
M949 211 221 225 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=29630 $D=0
M950 226 16 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=25000 $D=0
M951 227 16 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=29630 $D=0
M952 228 16 224 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=25000 $D=0
M953 229 16 225 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=29630 $D=0
M954 222 226 228 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=25000 $D=0
M955 223 227 229 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=29630 $D=0
M956 9 17 230 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=25000 $D=0
M957 9 17 231 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=29630 $D=0
M958 232 18 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=25000 $D=0
M959 233 18 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=29630 $D=0
M960 234 230 228 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=25000 $D=0
M961 235 231 229 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=29630 $D=0
M962 9 234 704 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=25000 $D=0
M963 9 235 705 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=29630 $D=0
M964 236 704 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=25000 $D=0
M965 237 705 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=29630 $D=0
M966 234 17 236 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=25000 $D=0
M967 235 17 237 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=29630 $D=0
M968 236 232 238 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=25000 $D=0
M969 237 233 239 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=29630 $D=0
M970 242 240 236 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=25000 $D=0
M971 243 241 237 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=29630 $D=0
M972 240 19 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=25000 $D=0
M973 241 19 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=29630 $D=0
M974 9 20 244 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=25000 $D=0
M975 9 20 245 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=29630 $D=0
M976 246 21 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=25000 $D=0
M977 247 21 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=29630 $D=0
M978 248 244 228 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=25000 $D=0
M979 249 245 229 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=29630 $D=0
M980 9 248 706 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=25000 $D=0
M981 9 249 707 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=29630 $D=0
M982 250 706 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=25000 $D=0
M983 251 707 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=29630 $D=0
M984 248 20 250 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=25000 $D=0
M985 249 20 251 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=29630 $D=0
M986 250 246 238 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=25000 $D=0
M987 251 247 239 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=29630 $D=0
M988 242 252 250 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=25000 $D=0
M989 243 253 251 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=29630 $D=0
M990 252 22 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=25000 $D=0
M991 253 22 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=29630 $D=0
M992 9 23 254 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=25000 $D=0
M993 9 23 255 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=29630 $D=0
M994 256 24 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=25000 $D=0
M995 257 24 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=29630 $D=0
M996 258 254 228 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=25000 $D=0
M997 259 255 229 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=29630 $D=0
M998 9 258 708 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=25000 $D=0
M999 9 259 709 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=29630 $D=0
M1000 260 708 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=25000 $D=0
M1001 261 709 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=29630 $D=0
M1002 258 23 260 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=25000 $D=0
M1003 259 23 261 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=29630 $D=0
M1004 260 256 238 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=25000 $D=0
M1005 261 257 239 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=29630 $D=0
M1006 242 262 260 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=25000 $D=0
M1007 243 263 261 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=29630 $D=0
M1008 262 25 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=25000 $D=0
M1009 263 25 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=29630 $D=0
M1010 9 26 264 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=25000 $D=0
M1011 9 26 265 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=29630 $D=0
M1012 266 27 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=25000 $D=0
M1013 267 27 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=29630 $D=0
M1014 268 264 228 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=25000 $D=0
M1015 269 265 229 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=29630 $D=0
M1016 9 268 710 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=25000 $D=0
M1017 9 269 711 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=29630 $D=0
M1018 270 710 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=25000 $D=0
M1019 271 711 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=29630 $D=0
M1020 268 26 270 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=25000 $D=0
M1021 269 26 271 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=29630 $D=0
M1022 270 266 238 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=25000 $D=0
M1023 271 267 239 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=29630 $D=0
M1024 242 272 270 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=25000 $D=0
M1025 243 273 271 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=29630 $D=0
M1026 272 28 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=25000 $D=0
M1027 273 28 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=29630 $D=0
M1028 9 29 274 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=25000 $D=0
M1029 9 29 275 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=29630 $D=0
M1030 276 30 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=25000 $D=0
M1031 277 30 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=29630 $D=0
M1032 278 274 228 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=25000 $D=0
M1033 279 275 229 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=29630 $D=0
M1034 9 278 712 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=25000 $D=0
M1035 9 279 713 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=29630 $D=0
M1036 280 712 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=25000 $D=0
M1037 281 713 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=29630 $D=0
M1038 278 29 280 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=25000 $D=0
M1039 279 29 281 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=29630 $D=0
M1040 280 276 238 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=25000 $D=0
M1041 281 277 239 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=29630 $D=0
M1042 242 282 280 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=25000 $D=0
M1043 243 283 281 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=29630 $D=0
M1044 282 31 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=25000 $D=0
M1045 283 31 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=29630 $D=0
M1046 9 32 284 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=25000 $D=0
M1047 9 32 285 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=29630 $D=0
M1048 286 33 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=25000 $D=0
M1049 287 33 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=29630 $D=0
M1050 288 284 228 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=25000 $D=0
M1051 289 285 229 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=29630 $D=0
M1052 9 288 714 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=25000 $D=0
M1053 9 289 715 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=29630 $D=0
M1054 290 714 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=25000 $D=0
M1055 291 715 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=29630 $D=0
M1056 288 32 290 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=25000 $D=0
M1057 289 32 291 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=29630 $D=0
M1058 290 286 238 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=25000 $D=0
M1059 291 287 239 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=29630 $D=0
M1060 242 292 290 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=25000 $D=0
M1061 243 293 291 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=29630 $D=0
M1062 292 34 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=25000 $D=0
M1063 293 34 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=29630 $D=0
M1064 9 35 294 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=25000 $D=0
M1065 9 35 295 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=29630 $D=0
M1066 296 36 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=25000 $D=0
M1067 297 36 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=29630 $D=0
M1068 298 294 228 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=25000 $D=0
M1069 299 295 229 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=29630 $D=0
M1070 9 298 716 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=25000 $D=0
M1071 9 299 717 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=29630 $D=0
M1072 300 716 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=25000 $D=0
M1073 301 717 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=29630 $D=0
M1074 298 35 300 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=25000 $D=0
M1075 299 35 301 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=29630 $D=0
M1076 300 296 238 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=25000 $D=0
M1077 301 297 239 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=29630 $D=0
M1078 242 302 300 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=25000 $D=0
M1079 243 303 301 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=29630 $D=0
M1080 302 37 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=25000 $D=0
M1081 303 37 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=29630 $D=0
M1082 9 38 304 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=25000 $D=0
M1083 9 38 305 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=29630 $D=0
M1084 306 39 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=25000 $D=0
M1085 307 39 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=29630 $D=0
M1086 308 304 228 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=25000 $D=0
M1087 309 305 229 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=29630 $D=0
M1088 9 308 718 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=25000 $D=0
M1089 9 309 719 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=29630 $D=0
M1090 310 718 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=25000 $D=0
M1091 311 719 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=29630 $D=0
M1092 308 38 310 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=25000 $D=0
M1093 309 38 311 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=29630 $D=0
M1094 310 306 238 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=25000 $D=0
M1095 311 307 239 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=29630 $D=0
M1096 242 312 310 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=25000 $D=0
M1097 243 313 311 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=29630 $D=0
M1098 312 40 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=25000 $D=0
M1099 313 40 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=29630 $D=0
M1100 9 41 314 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=25000 $D=0
M1101 9 41 315 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=29630 $D=0
M1102 316 42 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=25000 $D=0
M1103 317 42 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=29630 $D=0
M1104 318 314 228 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=25000 $D=0
M1105 319 315 229 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=29630 $D=0
M1106 9 318 720 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=25000 $D=0
M1107 9 319 721 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=29630 $D=0
M1108 320 720 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=25000 $D=0
M1109 321 721 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=29630 $D=0
M1110 318 41 320 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=25000 $D=0
M1111 319 41 321 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=29630 $D=0
M1112 320 316 238 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=25000 $D=0
M1113 321 317 239 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=29630 $D=0
M1114 242 322 320 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=25000 $D=0
M1115 243 323 321 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=29630 $D=0
M1116 322 43 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=25000 $D=0
M1117 323 43 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=29630 $D=0
M1118 9 44 324 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=25000 $D=0
M1119 9 44 325 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=29630 $D=0
M1120 326 45 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=25000 $D=0
M1121 327 45 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=29630 $D=0
M1122 328 324 228 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=25000 $D=0
M1123 329 325 229 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=29630 $D=0
M1124 9 328 722 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=25000 $D=0
M1125 9 329 723 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=29630 $D=0
M1126 330 722 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=25000 $D=0
M1127 331 723 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=29630 $D=0
M1128 328 44 330 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=25000 $D=0
M1129 329 44 331 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=29630 $D=0
M1130 330 326 238 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=25000 $D=0
M1131 331 327 239 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=29630 $D=0
M1132 242 332 330 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=25000 $D=0
M1133 243 333 331 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=29630 $D=0
M1134 332 46 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=25000 $D=0
M1135 333 46 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=29630 $D=0
M1136 9 47 334 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=25000 $D=0
M1137 9 47 335 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=29630 $D=0
M1138 336 48 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=25000 $D=0
M1139 337 48 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=29630 $D=0
M1140 338 334 228 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=25000 $D=0
M1141 339 335 229 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=29630 $D=0
M1142 9 338 724 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=25000 $D=0
M1143 9 339 725 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=29630 $D=0
M1144 340 724 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=25000 $D=0
M1145 341 725 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=29630 $D=0
M1146 338 47 340 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=25000 $D=0
M1147 339 47 341 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=29630 $D=0
M1148 340 336 238 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=25000 $D=0
M1149 341 337 239 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=29630 $D=0
M1150 242 342 340 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=25000 $D=0
M1151 243 343 341 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=29630 $D=0
M1152 342 49 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=25000 $D=0
M1153 343 49 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=29630 $D=0
M1154 9 50 344 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=25000 $D=0
M1155 9 50 345 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=29630 $D=0
M1156 346 51 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=25000 $D=0
M1157 347 51 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=29630 $D=0
M1158 348 344 228 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=25000 $D=0
M1159 349 345 229 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=29630 $D=0
M1160 9 348 726 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=25000 $D=0
M1161 9 349 727 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=29630 $D=0
M1162 350 726 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=25000 $D=0
M1163 351 727 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=29630 $D=0
M1164 348 50 350 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=25000 $D=0
M1165 349 50 351 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=29630 $D=0
M1166 350 346 238 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=25000 $D=0
M1167 351 347 239 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=29630 $D=0
M1168 242 352 350 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=25000 $D=0
M1169 243 353 351 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=29630 $D=0
M1170 352 52 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=25000 $D=0
M1171 353 52 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=29630 $D=0
M1172 9 53 354 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=25000 $D=0
M1173 9 53 355 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=29630 $D=0
M1174 356 54 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=25000 $D=0
M1175 357 54 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=29630 $D=0
M1176 358 354 228 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=25000 $D=0
M1177 359 355 229 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=29630 $D=0
M1178 9 358 728 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=25000 $D=0
M1179 9 359 729 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=29630 $D=0
M1180 360 728 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=25000 $D=0
M1181 361 729 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=29630 $D=0
M1182 358 53 360 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=25000 $D=0
M1183 359 53 361 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=29630 $D=0
M1184 360 356 238 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=25000 $D=0
M1185 361 357 239 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=29630 $D=0
M1186 242 362 360 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=25000 $D=0
M1187 243 363 361 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=29630 $D=0
M1188 362 55 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=25000 $D=0
M1189 363 55 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=29630 $D=0
M1190 9 56 364 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=25000 $D=0
M1191 9 56 365 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=29630 $D=0
M1192 366 57 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=25000 $D=0
M1193 367 57 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=29630 $D=0
M1194 368 364 228 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=25000 $D=0
M1195 369 365 229 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=29630 $D=0
M1196 9 368 730 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=25000 $D=0
M1197 9 369 731 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=29630 $D=0
M1198 370 730 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=25000 $D=0
M1199 371 731 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=29630 $D=0
M1200 368 56 370 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=25000 $D=0
M1201 369 56 371 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=29630 $D=0
M1202 370 366 238 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=25000 $D=0
M1203 371 367 239 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=29630 $D=0
M1204 242 372 370 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=25000 $D=0
M1205 243 373 371 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=29630 $D=0
M1206 372 58 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=25000 $D=0
M1207 373 58 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=29630 $D=0
M1208 9 59 374 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=25000 $D=0
M1209 9 59 375 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=29630 $D=0
M1210 376 60 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=25000 $D=0
M1211 377 60 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=29630 $D=0
M1212 378 374 228 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=25000 $D=0
M1213 379 375 229 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=29630 $D=0
M1214 9 378 732 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=25000 $D=0
M1215 9 379 733 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=29630 $D=0
M1216 380 732 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=25000 $D=0
M1217 381 733 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=29630 $D=0
M1218 378 59 380 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=25000 $D=0
M1219 379 59 381 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=29630 $D=0
M1220 380 376 238 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=25000 $D=0
M1221 381 377 239 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=29630 $D=0
M1222 242 382 380 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=25000 $D=0
M1223 243 383 381 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=29630 $D=0
M1224 382 61 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=25000 $D=0
M1225 383 61 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=29630 $D=0
M1226 9 62 384 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=25000 $D=0
M1227 9 62 385 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=29630 $D=0
M1228 386 63 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=25000 $D=0
M1229 387 63 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=29630 $D=0
M1230 388 384 228 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=25000 $D=0
M1231 389 385 229 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=29630 $D=0
M1232 9 388 734 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=25000 $D=0
M1233 9 389 735 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=29630 $D=0
M1234 390 734 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=25000 $D=0
M1235 391 735 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=29630 $D=0
M1236 388 62 390 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=25000 $D=0
M1237 389 62 391 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=29630 $D=0
M1238 390 386 238 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=25000 $D=0
M1239 391 387 239 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=29630 $D=0
M1240 242 392 390 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=25000 $D=0
M1241 243 393 391 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=29630 $D=0
M1242 392 64 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=25000 $D=0
M1243 393 64 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=29630 $D=0
M1244 9 65 394 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=25000 $D=0
M1245 9 65 395 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=29630 $D=0
M1246 396 66 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=25000 $D=0
M1247 397 66 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=29630 $D=0
M1248 398 394 228 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=25000 $D=0
M1249 399 395 229 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=29630 $D=0
M1250 9 398 736 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=25000 $D=0
M1251 9 399 737 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=29630 $D=0
M1252 400 736 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=25000 $D=0
M1253 401 737 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=29630 $D=0
M1254 398 65 400 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=25000 $D=0
M1255 399 65 401 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=29630 $D=0
M1256 400 396 238 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=25000 $D=0
M1257 401 397 239 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=29630 $D=0
M1258 242 402 400 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=25000 $D=0
M1259 243 403 401 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=29630 $D=0
M1260 402 67 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=25000 $D=0
M1261 403 67 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=29630 $D=0
M1262 9 68 404 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=25000 $D=0
M1263 9 68 405 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=29630 $D=0
M1264 406 69 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=25000 $D=0
M1265 407 69 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=29630 $D=0
M1266 408 404 228 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=25000 $D=0
M1267 409 405 229 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=29630 $D=0
M1268 9 408 738 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=25000 $D=0
M1269 9 409 739 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=29630 $D=0
M1270 410 738 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=25000 $D=0
M1271 411 739 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=29630 $D=0
M1272 408 68 410 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=25000 $D=0
M1273 409 68 411 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=29630 $D=0
M1274 410 406 238 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=25000 $D=0
M1275 411 407 239 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=29630 $D=0
M1276 242 412 410 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=25000 $D=0
M1277 243 413 411 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=29630 $D=0
M1278 412 70 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=25000 $D=0
M1279 413 70 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=29630 $D=0
M1280 9 71 414 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=25000 $D=0
M1281 9 71 415 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=29630 $D=0
M1282 416 72 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=25000 $D=0
M1283 417 72 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=29630 $D=0
M1284 418 414 228 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=25000 $D=0
M1285 419 415 229 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=29630 $D=0
M1286 9 418 740 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=25000 $D=0
M1287 9 419 741 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=29630 $D=0
M1288 420 740 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=25000 $D=0
M1289 421 741 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=29630 $D=0
M1290 418 71 420 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=25000 $D=0
M1291 419 71 421 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=29630 $D=0
M1292 420 416 238 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=25000 $D=0
M1293 421 417 239 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=29630 $D=0
M1294 242 422 420 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=25000 $D=0
M1295 243 423 421 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=29630 $D=0
M1296 422 73 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=25000 $D=0
M1297 423 73 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=29630 $D=0
M1298 9 74 424 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=25000 $D=0
M1299 9 74 425 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=29630 $D=0
M1300 426 75 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=25000 $D=0
M1301 427 75 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=29630 $D=0
M1302 428 424 228 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=25000 $D=0
M1303 429 425 229 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=29630 $D=0
M1304 9 428 742 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=25000 $D=0
M1305 9 429 743 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=29630 $D=0
M1306 430 742 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=25000 $D=0
M1307 431 743 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=29630 $D=0
M1308 428 74 430 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=25000 $D=0
M1309 429 74 431 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=29630 $D=0
M1310 430 426 238 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=25000 $D=0
M1311 431 427 239 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=29630 $D=0
M1312 242 432 430 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=25000 $D=0
M1313 243 433 431 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=29630 $D=0
M1314 432 76 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=25000 $D=0
M1315 433 76 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=29630 $D=0
M1316 9 77 434 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=25000 $D=0
M1317 9 77 435 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=29630 $D=0
M1318 436 78 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=25000 $D=0
M1319 437 78 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=29630 $D=0
M1320 438 434 228 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=25000 $D=0
M1321 439 435 229 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=29630 $D=0
M1322 9 438 744 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=25000 $D=0
M1323 9 439 745 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=29630 $D=0
M1324 440 744 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=25000 $D=0
M1325 441 745 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=29630 $D=0
M1326 438 77 440 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=25000 $D=0
M1327 439 77 441 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=29630 $D=0
M1328 440 436 238 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=25000 $D=0
M1329 441 437 239 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=29630 $D=0
M1330 242 442 440 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=25000 $D=0
M1331 243 443 441 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=29630 $D=0
M1332 442 79 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=25000 $D=0
M1333 443 79 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=29630 $D=0
M1334 9 80 444 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=25000 $D=0
M1335 9 80 445 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=29630 $D=0
M1336 446 81 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=25000 $D=0
M1337 447 81 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=29630 $D=0
M1338 448 444 228 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=25000 $D=0
M1339 449 445 229 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=29630 $D=0
M1340 9 448 746 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=25000 $D=0
M1341 9 449 747 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=29630 $D=0
M1342 450 746 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=25000 $D=0
M1343 451 747 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=29630 $D=0
M1344 448 80 450 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=25000 $D=0
M1345 449 80 451 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=29630 $D=0
M1346 450 446 238 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=25000 $D=0
M1347 451 447 239 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=29630 $D=0
M1348 242 452 450 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=25000 $D=0
M1349 243 453 451 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=29630 $D=0
M1350 452 82 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=25000 $D=0
M1351 453 82 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=29630 $D=0
M1352 9 83 454 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=25000 $D=0
M1353 9 83 455 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=29630 $D=0
M1354 456 84 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=25000 $D=0
M1355 457 84 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=29630 $D=0
M1356 458 454 228 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=25000 $D=0
M1357 459 455 229 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=29630 $D=0
M1358 9 458 748 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=25000 $D=0
M1359 9 459 749 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=29630 $D=0
M1360 460 748 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=25000 $D=0
M1361 461 749 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=29630 $D=0
M1362 458 83 460 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=25000 $D=0
M1363 459 83 461 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=29630 $D=0
M1364 460 456 238 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=25000 $D=0
M1365 461 457 239 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=29630 $D=0
M1366 242 462 460 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=25000 $D=0
M1367 243 463 461 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=29630 $D=0
M1368 462 85 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=25000 $D=0
M1369 463 85 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=29630 $D=0
M1370 9 86 464 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=25000 $D=0
M1371 9 86 465 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=29630 $D=0
M1372 466 87 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=25000 $D=0
M1373 467 87 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=29630 $D=0
M1374 468 464 228 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=25000 $D=0
M1375 469 465 229 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=29630 $D=0
M1376 9 468 750 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=25000 $D=0
M1377 9 469 751 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=29630 $D=0
M1378 470 750 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=25000 $D=0
M1379 471 751 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=29630 $D=0
M1380 468 86 470 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=25000 $D=0
M1381 469 86 471 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=29630 $D=0
M1382 470 466 238 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=25000 $D=0
M1383 471 467 239 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=29630 $D=0
M1384 242 472 470 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=25000 $D=0
M1385 243 473 471 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=29630 $D=0
M1386 472 88 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=25000 $D=0
M1387 473 88 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=29630 $D=0
M1388 9 89 474 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=25000 $D=0
M1389 9 89 475 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=29630 $D=0
M1390 476 90 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=25000 $D=0
M1391 477 90 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=29630 $D=0
M1392 478 474 228 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=25000 $D=0
M1393 479 475 229 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=29630 $D=0
M1394 9 478 752 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=25000 $D=0
M1395 9 479 753 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=29630 $D=0
M1396 480 752 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=25000 $D=0
M1397 481 753 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=29630 $D=0
M1398 478 89 480 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=25000 $D=0
M1399 479 89 481 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=29630 $D=0
M1400 480 476 238 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=25000 $D=0
M1401 481 477 239 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=29630 $D=0
M1402 242 482 480 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=25000 $D=0
M1403 243 483 481 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=29630 $D=0
M1404 482 91 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=25000 $D=0
M1405 483 91 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=29630 $D=0
M1406 9 92 484 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=25000 $D=0
M1407 9 92 485 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=29630 $D=0
M1408 486 93 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=25000 $D=0
M1409 487 93 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=29630 $D=0
M1410 488 484 228 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=25000 $D=0
M1411 489 485 229 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=29630 $D=0
M1412 9 488 754 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=25000 $D=0
M1413 9 489 755 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=29630 $D=0
M1414 490 754 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=25000 $D=0
M1415 491 755 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=29630 $D=0
M1416 488 92 490 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=25000 $D=0
M1417 489 92 491 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=29630 $D=0
M1418 490 486 238 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=25000 $D=0
M1419 491 487 239 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=29630 $D=0
M1420 242 492 490 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=25000 $D=0
M1421 243 493 491 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=29630 $D=0
M1422 492 94 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=25000 $D=0
M1423 493 94 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=29630 $D=0
M1424 9 95 494 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=25000 $D=0
M1425 9 95 495 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=29630 $D=0
M1426 496 96 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=25000 $D=0
M1427 497 96 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=29630 $D=0
M1428 498 494 228 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=25000 $D=0
M1429 499 495 229 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=29630 $D=0
M1430 9 498 756 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=25000 $D=0
M1431 9 499 757 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=29630 $D=0
M1432 500 756 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=25000 $D=0
M1433 501 757 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=29630 $D=0
M1434 498 95 500 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=25000 $D=0
M1435 499 95 501 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=29630 $D=0
M1436 500 496 238 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=25000 $D=0
M1437 501 497 239 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=29630 $D=0
M1438 242 502 500 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=25000 $D=0
M1439 243 503 501 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=29630 $D=0
M1440 502 97 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=25000 $D=0
M1441 503 97 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=29630 $D=0
M1442 9 98 504 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=25000 $D=0
M1443 9 98 505 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=29630 $D=0
M1444 506 99 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=25000 $D=0
M1445 507 99 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=29630 $D=0
M1446 508 504 228 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=25000 $D=0
M1447 509 505 229 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=29630 $D=0
M1448 9 508 758 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=25000 $D=0
M1449 9 509 759 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=29630 $D=0
M1450 510 758 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=25000 $D=0
M1451 511 759 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=29630 $D=0
M1452 508 98 510 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=25000 $D=0
M1453 509 98 511 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=29630 $D=0
M1454 510 506 238 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=25000 $D=0
M1455 511 507 239 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=29630 $D=0
M1456 242 512 510 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=25000 $D=0
M1457 243 513 511 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=29630 $D=0
M1458 512 100 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=25000 $D=0
M1459 513 100 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=29630 $D=0
M1460 9 101 514 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=25000 $D=0
M1461 9 101 515 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=29630 $D=0
M1462 516 102 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=25000 $D=0
M1463 517 102 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=29630 $D=0
M1464 518 514 228 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=25000 $D=0
M1465 519 515 229 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=29630 $D=0
M1466 9 518 760 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=25000 $D=0
M1467 9 519 761 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=29630 $D=0
M1468 520 760 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=25000 $D=0
M1469 521 761 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=29630 $D=0
M1470 518 101 520 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=25000 $D=0
M1471 519 101 521 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=29630 $D=0
M1472 520 516 238 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=25000 $D=0
M1473 521 517 239 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=29630 $D=0
M1474 242 522 520 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=25000 $D=0
M1475 243 523 521 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=29630 $D=0
M1476 522 103 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=25000 $D=0
M1477 523 103 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=29630 $D=0
M1478 9 104 524 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=25000 $D=0
M1479 9 104 525 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=29630 $D=0
M1480 526 105 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=25000 $D=0
M1481 527 105 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=29630 $D=0
M1482 528 524 228 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=25000 $D=0
M1483 529 525 229 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=29630 $D=0
M1484 9 528 762 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=25000 $D=0
M1485 9 529 763 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=29630 $D=0
M1486 530 762 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=25000 $D=0
M1487 531 763 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=29630 $D=0
M1488 528 104 530 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=25000 $D=0
M1489 529 104 531 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=29630 $D=0
M1490 530 526 238 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=25000 $D=0
M1491 531 527 239 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=29630 $D=0
M1492 242 532 530 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=25000 $D=0
M1493 243 533 531 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=29630 $D=0
M1494 532 107 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=25000 $D=0
M1495 533 107 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=29630 $D=0
M1496 9 108 534 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=25000 $D=0
M1497 9 108 535 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=29630 $D=0
M1498 536 109 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=25000 $D=0
M1499 537 109 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=29630 $D=0
M1500 538 534 228 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=25000 $D=0
M1501 539 535 229 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=29630 $D=0
M1502 9 538 764 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=25000 $D=0
M1503 9 539 765 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=29630 $D=0
M1504 540 764 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=25000 $D=0
M1505 541 765 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=29630 $D=0
M1506 538 108 540 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=25000 $D=0
M1507 539 108 541 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=29630 $D=0
M1508 540 536 238 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=25000 $D=0
M1509 541 537 239 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=29630 $D=0
M1510 242 542 540 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=25000 $D=0
M1511 243 543 541 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=29630 $D=0
M1512 542 111 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=25000 $D=0
M1513 543 111 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=29630 $D=0
M1514 9 112 544 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=25000 $D=0
M1515 9 112 545 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=29630 $D=0
M1516 546 113 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=25000 $D=0
M1517 547 113 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=29630 $D=0
M1518 6 546 238 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=25000 $D=0
M1519 6 547 239 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=29630 $D=0
M1520 242 544 6 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=25000 $D=0
M1521 243 545 6 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=29630 $D=0
M1522 9 550 548 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=25000 $D=0
M1523 9 551 549 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=29630 $D=0
M1524 550 115 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=25000 $D=0
M1525 551 115 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=29630 $D=0
M1526 766 238 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=25000 $D=0
M1527 767 239 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=29630 $D=0
M1528 552 550 766 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=25000 $D=0
M1529 553 551 767 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=29630 $D=0
M1530 9 552 554 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=25000 $D=0
M1531 9 553 555 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=29630 $D=0
M1532 768 554 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=25000 $D=0
M1533 769 555 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=29630 $D=0
M1534 552 548 768 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=25000 $D=0
M1535 553 549 769 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=29630 $D=0
M1536 9 558 556 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=25000 $D=0
M1537 9 559 557 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=29630 $D=0
M1538 558 115 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=25000 $D=0
M1539 559 115 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=29630 $D=0
M1540 770 242 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=25000 $D=0
M1541 771 243 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=29630 $D=0
M1542 560 558 770 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=25000 $D=0
M1543 561 559 771 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=29630 $D=0
M1544 9 560 117 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=25000 $D=0
M1545 9 561 118 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=29630 $D=0
M1546 772 117 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=25000 $D=0
M1547 773 118 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=29630 $D=0
M1548 560 556 772 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=25000 $D=0
M1549 561 557 773 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=29630 $D=0
M1550 562 119 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=25000 $D=0
M1551 563 119 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=29630 $D=0
M1552 564 119 554 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=25000 $D=0
M1553 565 119 555 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=29630 $D=0
M1554 120 562 564 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=25000 $D=0
M1555 121 563 565 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=29630 $D=0
M1556 566 122 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=25000 $D=0
M1557 567 122 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=29630 $D=0
M1558 568 122 117 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=25000 $D=0
M1559 569 122 118 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=29630 $D=0
M1560 774 566 568 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=25000 $D=0
M1561 775 567 569 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=29630 $D=0
M1562 9 117 774 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=25000 $D=0
M1563 9 118 775 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=29630 $D=0
M1564 570 123 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=25000 $D=0
M1565 571 123 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=29630 $D=0
M1566 572 123 568 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=25000 $D=0
M1567 573 123 569 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=29630 $D=0
M1568 11 570 572 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=25000 $D=0
M1569 12 571 573 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=29630 $D=0
M1570 575 574 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=25000 $D=0
M1571 576 124 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=29630 $D=0
M1572 9 579 577 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=25000 $D=0
M1573 9 580 578 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=29630 $D=0
M1574 581 564 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=25000 $D=0
M1575 582 565 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=29630 $D=0
M1576 579 564 574 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=25000 $D=0
M1577 580 565 124 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=29630 $D=0
M1578 575 581 579 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=25000 $D=0
M1579 576 582 580 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=29630 $D=0
M1580 583 577 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=25000 $D=0
M1581 584 578 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=29630 $D=0
M1582 125 577 572 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=25000 $D=0
M1583 574 578 573 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=29630 $D=0
M1584 564 583 125 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=25000 $D=0
M1585 565 584 574 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=29630 $D=0
M1586 585 125 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=25000 $D=0
M1587 586 574 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=29630 $D=0
M1588 587 577 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=25000 $D=0
M1589 588 578 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=29630 $D=0
M1590 589 577 585 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=25000 $D=0
M1591 590 578 586 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=29630 $D=0
M1592 572 587 589 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=25000 $D=0
M1593 573 588 590 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=29630 $D=0
M1594 786 564 9 9 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=24640 $D=0
M1595 787 565 9 9 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=29270 $D=0
M1596 591 572 786 9 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=24640 $D=0
M1597 592 573 787 9 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=29270 $D=0
M1598 593 589 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=25000 $D=0
M1599 594 590 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=29630 $D=0
M1600 595 564 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=25000 $D=0
M1601 596 565 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=29630 $D=0
M1602 9 572 595 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=25000 $D=0
M1603 9 573 596 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=29630 $D=0
M1604 597 564 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=25000 $D=0
M1605 598 565 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=29630 $D=0
M1606 9 572 597 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=25000 $D=0
M1607 9 573 598 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=29630 $D=0
M1608 788 564 9 9 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=24820 $D=0
M1609 789 565 9 9 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=29450 $D=0
M1610 601 572 788 9 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=24820 $D=0
M1611 602 573 789 9 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=29450 $D=0
M1612 9 597 601 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=25000 $D=0
M1613 9 598 602 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=29630 $D=0
M1614 603 128 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=25000 $D=0
M1615 604 128 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=29630 $D=0
M1616 605 128 591 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=25000 $D=0
M1617 606 128 592 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=29630 $D=0
M1618 595 603 605 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=25000 $D=0
M1619 596 604 606 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=29630 $D=0
M1620 607 128 593 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=25000 $D=0
M1621 608 128 594 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=29630 $D=0
M1622 601 603 607 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=25000 $D=0
M1623 602 604 608 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=29630 $D=0
M1624 609 129 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=25000 $D=0
M1625 610 129 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=29630 $D=0
M1626 611 129 607 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=25000 $D=0
M1627 612 129 608 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=29630 $D=0
M1628 605 609 611 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=25000 $D=0
M1629 606 610 612 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=29630 $D=0
M1630 13 611 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=25000 $D=0
M1631 14 612 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=29630 $D=0
M1632 613 130 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=25000 $D=0
M1633 614 130 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=29630 $D=0
M1634 615 130 131 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=25000 $D=0
M1635 616 130 132 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=29630 $D=0
M1636 133 613 615 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=25000 $D=0
M1637 134 614 616 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=29630 $D=0
M1638 617 130 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=25000 $D=0
M1639 618 130 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=29630 $D=0
M1640 619 130 135 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=25000 $D=0
M1641 620 130 136 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=29630 $D=0
M1642 137 617 619 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=25000 $D=0
M1643 138 618 620 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=29630 $D=0
M1644 621 130 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=25000 $D=0
M1645 622 130 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=29630 $D=0
M1646 623 130 127 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=25000 $D=0
M1647 624 130 126 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=29630 $D=0
M1648 139 621 623 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=25000 $D=0
M1649 140 622 624 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=29630 $D=0
M1650 625 130 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=25000 $D=0
M1651 626 130 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=29630 $D=0
M1652 627 130 142 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=25000 $D=0
M1653 628 130 143 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=29630 $D=0
M1654 144 625 627 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=25000 $D=0
M1655 144 626 628 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=29630 $D=0
M1656 629 130 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=25000 $D=0
M1657 630 130 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=29630 $D=0
M1658 631 130 145 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=25000 $D=0
M1659 632 130 146 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=29630 $D=0
M1660 144 629 631 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=25000 $D=0
M1661 144 630 632 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=29630 $D=0
M1662 9 564 776 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=25000 $D=0
M1663 9 565 777 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=29630 $D=0
M1664 134 776 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=25000 $D=0
M1665 131 777 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=29630 $D=0
M1666 633 147 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=25000 $D=0
M1667 634 147 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=29630 $D=0
M1668 148 147 134 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=25000 $D=0
M1669 149 147 131 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=29630 $D=0
M1670 615 633 148 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=25000 $D=0
M1671 616 634 149 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=29630 $D=0
M1672 635 150 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=25000 $D=0
M1673 636 150 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=29630 $D=0
M1674 151 150 148 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=25000 $D=0
M1675 106 150 149 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=29630 $D=0
M1676 619 635 151 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=25000 $D=0
M1677 620 636 106 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=29630 $D=0
M1678 637 152 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=25000 $D=0
M1679 638 152 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=29630 $D=0
M1680 153 152 151 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=25000 $D=0
M1681 114 152 106 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=29630 $D=0
M1682 623 637 153 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=25000 $D=0
M1683 624 638 114 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=29630 $D=0
M1684 639 154 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=25000 $D=0
M1685 640 154 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=29630 $D=0
M1686 155 154 153 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=25000 $D=0
M1687 156 154 114 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=29630 $D=0
M1688 627 639 155 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=25000 $D=0
M1689 628 640 156 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=29630 $D=0
M1690 641 157 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=25000 $D=0
M1691 642 157 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=29630 $D=0
M1692 214 157 155 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=25000 $D=0
M1693 215 157 156 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=29630 $D=0
M1694 631 641 214 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=25000 $D=0
M1695 632 642 215 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=29630 $D=0
M1696 643 158 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=25000 $D=0
M1697 644 158 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=29630 $D=0
M1698 645 158 117 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=25000 $D=0
M1699 646 158 118 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=29630 $D=0
M1700 11 643 645 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=25000 $D=0
M1701 12 644 646 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=29630 $D=0
M1702 647 554 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=25000 $D=0
M1703 648 555 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=29630 $D=0
M1704 9 645 647 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=25000 $D=0
M1705 9 646 648 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=29630 $D=0
M1706 790 554 9 9 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=24820 $D=0
M1707 791 555 9 9 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=29450 $D=0
M1708 651 645 790 9 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=24820 $D=0
M1709 652 646 791 9 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=29450 $D=0
M1710 9 647 651 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=25000 $D=0
M1711 9 648 652 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=29630 $D=0
M1712 778 159 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=25000 $D=0
M1713 779 653 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=29630 $D=0
M1714 9 651 778 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=25000 $D=0
M1715 9 652 779 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=29630 $D=0
M1716 653 778 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=25000 $D=0
M1717 160 779 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=29630 $D=0
M1718 792 554 9 9 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=24640 $D=0
M1719 793 555 9 9 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=29270 $D=0
M1720 654 656 792 9 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=24640 $D=0
M1721 655 657 793 9 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=29270 $D=0
M1722 656 645 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=25000 $D=0
M1723 657 646 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=29630 $D=0
M1724 658 654 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=25000 $D=0
M1725 659 655 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=29630 $D=0
M1726 9 159 658 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=25000 $D=0
M1727 9 653 659 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=29630 $D=0
M1728 661 161 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=25000 $D=0
M1729 662 660 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=29630 $D=0
M1730 660 658 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=25000 $D=0
M1731 162 659 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=29630 $D=0
M1732 9 661 660 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=25000 $D=0
M1733 9 662 162 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=29630 $D=0
M1734 664 663 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=25000 $D=0
M1735 665 163 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=29630 $D=0
M1736 9 668 666 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=25000 $D=0
M1737 9 669 667 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=29630 $D=0
M1738 670 120 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=25000 $D=0
M1739 671 121 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=29630 $D=0
M1740 668 120 663 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=25000 $D=0
M1741 669 121 163 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=29630 $D=0
M1742 664 670 668 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=25000 $D=0
M1743 665 671 669 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=29630 $D=0
M1744 672 666 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=25000 $D=0
M1745 673 667 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=29630 $D=0
M1746 164 666 6 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=25000 $D=0
M1747 663 667 6 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=29630 $D=0
M1748 120 672 164 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=25000 $D=0
M1749 121 673 663 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=29630 $D=0
M1750 674 164 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=25000 $D=0
M1751 675 663 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=29630 $D=0
M1752 676 666 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=25000 $D=0
M1753 677 667 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=29630 $D=0
M1754 216 666 674 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=25000 $D=0
M1755 217 667 675 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=29630 $D=0
M1756 6 676 216 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=25000 $D=0
M1757 6 677 217 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=29630 $D=0
M1758 678 165 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=25000 $D=0
M1759 679 165 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=29630 $D=0
M1760 680 165 216 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=25000 $D=0
M1761 681 165 217 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=29630 $D=0
M1762 13 678 680 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=25000 $D=0
M1763 14 679 681 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=29630 $D=0
M1764 682 166 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=25000 $D=0
M1765 683 166 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=29630 $D=0
M1766 684 166 680 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=25000 $D=0
M1767 685 166 681 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=29630 $D=0
M1768 6 682 684 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=25000 $D=0
M1769 6 683 685 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=29630 $D=0
M1770 686 115 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=25000 $D=0
M1771 687 115 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=29630 $D=0
M1772 9 686 688 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=25000 $D=0
M1773 9 687 689 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=29630 $D=0
M1774 690 115 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=25000 $D=0
M1775 691 115 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=29630 $D=0
M1776 692 688 684 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=25000 $D=0
M1777 693 689 685 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=29630 $D=0
M1778 9 692 780 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=25000 $D=0
M1779 9 693 781 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=29630 $D=0
M1780 694 780 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=25000 $D=0
M1781 695 781 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=29630 $D=0
M1782 692 686 694 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=25000 $D=0
M1783 693 687 695 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=29630 $D=0
M1784 696 690 694 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=25000 $D=0
M1785 697 691 695 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=29630 $D=0
M1786 9 700 698 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=25000 $D=0
M1787 9 701 699 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=29630 $D=0
M1788 700 115 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=25000 $D=0
M1789 701 115 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=29630 $D=0
M1790 782 696 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=25000 $D=0
M1791 783 697 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=29630 $D=0
M1792 702 700 782 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=25000 $D=0
M1793 703 701 783 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=29630 $D=0
M1794 9 702 120 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=25000 $D=0
M1795 9 703 121 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=29630 $D=0
M1796 784 120 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=25000 $D=0
M1797 785 121 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=29630 $D=0
M1798 702 698 784 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=25000 $D=0
M1799 703 699 785 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=29630 $D=0
.ENDS
***************************************
.SUBCKT ICV_40 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 109 110 111 113 114 115 116 117 118 119 120 121 122
+ 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 142 143
+ 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162 163
+ 164 165
** N=796 EP=162 IP=1514 FDC=1800
M0 181 1 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=14490 $D=1
M1 182 1 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=19120 $D=1
M2 183 181 2 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=14490 $D=1
M3 184 182 3 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=19120 $D=1
M4 6 1 183 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=14490 $D=1
M5 6 1 184 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=19120 $D=1
M6 185 181 4 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=14490 $D=1
M7 186 182 4 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=19120 $D=1
M8 5 1 185 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=14490 $D=1
M9 5 1 186 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=19120 $D=1
M10 187 181 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=14490 $D=1
M11 188 182 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=19120 $D=1
M12 6 1 187 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=14490 $D=1
M13 6 1 188 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=19120 $D=1
M14 191 189 187 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=14490 $D=1
M15 192 190 188 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=19120 $D=1
M16 189 7 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=14490 $D=1
M17 190 7 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=19120 $D=1
M18 193 189 185 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=14490 $D=1
M19 194 190 186 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=19120 $D=1
M20 183 7 193 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=14490 $D=1
M21 184 7 194 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=19120 $D=1
M22 195 8 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=14490 $D=1
M23 196 8 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=19120 $D=1
M24 197 195 193 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=14490 $D=1
M25 198 196 194 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=19120 $D=1
M26 191 8 197 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=14490 $D=1
M27 192 8 198 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=19120 $D=1
M28 199 10 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=14490 $D=1
M29 200 10 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=19120 $D=1
M30 201 199 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=14490 $D=1
M31 202 200 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=19120 $D=1
M32 11 10 201 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=14490 $D=1
M33 12 10 202 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=19120 $D=1
M34 203 199 13 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=14490 $D=1
M35 204 200 14 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=19120 $D=1
M36 205 10 203 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=14490 $D=1
M37 206 10 204 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=19120 $D=1
M38 209 199 207 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=14490 $D=1
M39 210 200 208 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=19120 $D=1
M40 197 10 209 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=14490 $D=1
M41 198 10 210 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=19120 $D=1
M42 213 211 209 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=14490 $D=1
M43 214 212 210 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=19120 $D=1
M44 211 15 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=14490 $D=1
M45 212 15 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=19120 $D=1
M46 215 211 203 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=14490 $D=1
M47 216 212 204 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=19120 $D=1
M48 201 15 215 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=14490 $D=1
M49 202 15 216 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=19120 $D=1
M50 217 16 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=14490 $D=1
M51 218 16 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=19120 $D=1
M52 219 217 215 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=14490 $D=1
M53 220 218 216 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=19120 $D=1
M54 213 16 219 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=14490 $D=1
M55 214 16 220 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=19120 $D=1
M56 6 17 221 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=14490 $D=1
M57 6 17 222 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=19120 $D=1
M58 223 18 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=14490 $D=1
M59 224 18 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=19120 $D=1
M60 225 17 219 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=14490 $D=1
M61 226 17 220 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=19120 $D=1
M62 6 225 695 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=14490 $D=1
M63 6 226 696 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=19120 $D=1
M64 227 695 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=14490 $D=1
M65 228 696 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=19120 $D=1
M66 225 221 227 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=14490 $D=1
M67 226 222 228 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=19120 $D=1
M68 227 18 229 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=14490 $D=1
M69 228 18 230 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=19120 $D=1
M70 233 19 227 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=14490 $D=1
M71 234 19 228 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=19120 $D=1
M72 231 19 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=14490 $D=1
M73 232 19 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=19120 $D=1
M74 6 20 235 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=14490 $D=1
M75 6 20 236 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=19120 $D=1
M76 237 21 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=14490 $D=1
M77 238 21 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=19120 $D=1
M78 239 20 219 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=14490 $D=1
M79 240 20 220 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=19120 $D=1
M80 6 239 697 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=14490 $D=1
M81 6 240 698 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=19120 $D=1
M82 241 697 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=14490 $D=1
M83 242 698 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=19120 $D=1
M84 239 235 241 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=14490 $D=1
M85 240 236 242 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=19120 $D=1
M86 241 21 229 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=14490 $D=1
M87 242 21 230 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=19120 $D=1
M88 233 22 241 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=14490 $D=1
M89 234 22 242 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=19120 $D=1
M90 243 22 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=14490 $D=1
M91 244 22 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=19120 $D=1
M92 6 23 245 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=14490 $D=1
M93 6 23 246 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=19120 $D=1
M94 247 24 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=14490 $D=1
M95 248 24 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=19120 $D=1
M96 249 23 219 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=14490 $D=1
M97 250 23 220 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=19120 $D=1
M98 6 249 699 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=14490 $D=1
M99 6 250 700 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=19120 $D=1
M100 251 699 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=14490 $D=1
M101 252 700 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=19120 $D=1
M102 249 245 251 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=14490 $D=1
M103 250 246 252 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=19120 $D=1
M104 251 24 229 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=14490 $D=1
M105 252 24 230 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=19120 $D=1
M106 233 25 251 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=14490 $D=1
M107 234 25 252 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=19120 $D=1
M108 253 25 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=14490 $D=1
M109 254 25 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=19120 $D=1
M110 6 26 255 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=14490 $D=1
M111 6 26 256 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=19120 $D=1
M112 257 27 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=14490 $D=1
M113 258 27 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=19120 $D=1
M114 259 26 219 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=14490 $D=1
M115 260 26 220 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=19120 $D=1
M116 6 259 701 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=14490 $D=1
M117 6 260 702 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=19120 $D=1
M118 261 701 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=14490 $D=1
M119 262 702 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=19120 $D=1
M120 259 255 261 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=14490 $D=1
M121 260 256 262 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=19120 $D=1
M122 261 27 229 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=14490 $D=1
M123 262 27 230 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=19120 $D=1
M124 233 28 261 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=14490 $D=1
M125 234 28 262 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=19120 $D=1
M126 263 28 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=14490 $D=1
M127 264 28 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=19120 $D=1
M128 6 29 265 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=14490 $D=1
M129 6 29 266 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=19120 $D=1
M130 267 30 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=14490 $D=1
M131 268 30 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=19120 $D=1
M132 269 29 219 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=14490 $D=1
M133 270 29 220 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=19120 $D=1
M134 6 269 703 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=14490 $D=1
M135 6 270 704 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=19120 $D=1
M136 271 703 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=14490 $D=1
M137 272 704 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=19120 $D=1
M138 269 265 271 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=14490 $D=1
M139 270 266 272 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=19120 $D=1
M140 271 30 229 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=14490 $D=1
M141 272 30 230 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=19120 $D=1
M142 233 31 271 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=14490 $D=1
M143 234 31 272 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=19120 $D=1
M144 273 31 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=14490 $D=1
M145 274 31 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=19120 $D=1
M146 6 32 275 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=14490 $D=1
M147 6 32 276 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=19120 $D=1
M148 277 33 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=14490 $D=1
M149 278 33 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=19120 $D=1
M150 279 32 219 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=14490 $D=1
M151 280 32 220 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=19120 $D=1
M152 6 279 705 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=14490 $D=1
M153 6 280 706 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=19120 $D=1
M154 281 705 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=14490 $D=1
M155 282 706 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=19120 $D=1
M156 279 275 281 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=14490 $D=1
M157 280 276 282 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=19120 $D=1
M158 281 33 229 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=14490 $D=1
M159 282 33 230 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=19120 $D=1
M160 233 34 281 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=14490 $D=1
M161 234 34 282 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=19120 $D=1
M162 283 34 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=14490 $D=1
M163 284 34 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=19120 $D=1
M164 6 35 285 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=14490 $D=1
M165 6 35 286 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=19120 $D=1
M166 287 36 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=14490 $D=1
M167 288 36 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=19120 $D=1
M168 289 35 219 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=14490 $D=1
M169 290 35 220 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=19120 $D=1
M170 6 289 707 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=14490 $D=1
M171 6 290 708 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=19120 $D=1
M172 291 707 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=14490 $D=1
M173 292 708 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=19120 $D=1
M174 289 285 291 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=14490 $D=1
M175 290 286 292 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=19120 $D=1
M176 291 36 229 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=14490 $D=1
M177 292 36 230 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=19120 $D=1
M178 233 37 291 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=14490 $D=1
M179 234 37 292 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=19120 $D=1
M180 293 37 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=14490 $D=1
M181 294 37 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=19120 $D=1
M182 6 38 295 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=14490 $D=1
M183 6 38 296 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=19120 $D=1
M184 297 39 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=14490 $D=1
M185 298 39 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=19120 $D=1
M186 299 38 219 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=14490 $D=1
M187 300 38 220 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=19120 $D=1
M188 6 299 709 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=14490 $D=1
M189 6 300 710 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=19120 $D=1
M190 301 709 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=14490 $D=1
M191 302 710 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=19120 $D=1
M192 299 295 301 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=14490 $D=1
M193 300 296 302 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=19120 $D=1
M194 301 39 229 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=14490 $D=1
M195 302 39 230 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=19120 $D=1
M196 233 40 301 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=14490 $D=1
M197 234 40 302 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=19120 $D=1
M198 303 40 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=14490 $D=1
M199 304 40 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=19120 $D=1
M200 6 41 305 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=14490 $D=1
M201 6 41 306 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=19120 $D=1
M202 307 42 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=14490 $D=1
M203 308 42 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=19120 $D=1
M204 309 41 219 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=14490 $D=1
M205 310 41 220 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=19120 $D=1
M206 6 309 711 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=14490 $D=1
M207 6 310 712 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=19120 $D=1
M208 311 711 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=14490 $D=1
M209 312 712 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=19120 $D=1
M210 309 305 311 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=14490 $D=1
M211 310 306 312 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=19120 $D=1
M212 311 42 229 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=14490 $D=1
M213 312 42 230 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=19120 $D=1
M214 233 43 311 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=14490 $D=1
M215 234 43 312 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=19120 $D=1
M216 313 43 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=14490 $D=1
M217 314 43 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=19120 $D=1
M218 6 44 315 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=14490 $D=1
M219 6 44 316 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=19120 $D=1
M220 317 45 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=14490 $D=1
M221 318 45 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=19120 $D=1
M222 319 44 219 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=14490 $D=1
M223 320 44 220 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=19120 $D=1
M224 6 319 713 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=14490 $D=1
M225 6 320 714 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=19120 $D=1
M226 321 713 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=14490 $D=1
M227 322 714 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=19120 $D=1
M228 319 315 321 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=14490 $D=1
M229 320 316 322 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=19120 $D=1
M230 321 45 229 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=14490 $D=1
M231 322 45 230 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=19120 $D=1
M232 233 46 321 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=14490 $D=1
M233 234 46 322 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=19120 $D=1
M234 323 46 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=14490 $D=1
M235 324 46 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=19120 $D=1
M236 6 47 325 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=14490 $D=1
M237 6 47 326 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=19120 $D=1
M238 327 48 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=14490 $D=1
M239 328 48 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=19120 $D=1
M240 329 47 219 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=14490 $D=1
M241 330 47 220 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=19120 $D=1
M242 6 329 715 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=14490 $D=1
M243 6 330 716 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=19120 $D=1
M244 331 715 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=14490 $D=1
M245 332 716 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=19120 $D=1
M246 329 325 331 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=14490 $D=1
M247 330 326 332 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=19120 $D=1
M248 331 48 229 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=14490 $D=1
M249 332 48 230 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=19120 $D=1
M250 233 49 331 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=14490 $D=1
M251 234 49 332 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=19120 $D=1
M252 333 49 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=14490 $D=1
M253 334 49 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=19120 $D=1
M254 6 50 335 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=14490 $D=1
M255 6 50 336 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=19120 $D=1
M256 337 51 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=14490 $D=1
M257 338 51 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=19120 $D=1
M258 339 50 219 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=14490 $D=1
M259 340 50 220 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=19120 $D=1
M260 6 339 717 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=14490 $D=1
M261 6 340 718 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=19120 $D=1
M262 341 717 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=14490 $D=1
M263 342 718 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=19120 $D=1
M264 339 335 341 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=14490 $D=1
M265 340 336 342 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=19120 $D=1
M266 341 51 229 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=14490 $D=1
M267 342 51 230 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=19120 $D=1
M268 233 52 341 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=14490 $D=1
M269 234 52 342 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=19120 $D=1
M270 343 52 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=14490 $D=1
M271 344 52 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=19120 $D=1
M272 6 53 345 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=14490 $D=1
M273 6 53 346 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=19120 $D=1
M274 347 54 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=14490 $D=1
M275 348 54 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=19120 $D=1
M276 349 53 219 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=14490 $D=1
M277 350 53 220 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=19120 $D=1
M278 6 349 719 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=14490 $D=1
M279 6 350 720 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=19120 $D=1
M280 351 719 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=14490 $D=1
M281 352 720 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=19120 $D=1
M282 349 345 351 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=14490 $D=1
M283 350 346 352 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=19120 $D=1
M284 351 54 229 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=14490 $D=1
M285 352 54 230 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=19120 $D=1
M286 233 55 351 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=14490 $D=1
M287 234 55 352 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=19120 $D=1
M288 353 55 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=14490 $D=1
M289 354 55 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=19120 $D=1
M290 6 56 355 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=14490 $D=1
M291 6 56 356 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=19120 $D=1
M292 357 57 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=14490 $D=1
M293 358 57 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=19120 $D=1
M294 359 56 219 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=14490 $D=1
M295 360 56 220 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=19120 $D=1
M296 6 359 721 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=14490 $D=1
M297 6 360 722 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=19120 $D=1
M298 361 721 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=14490 $D=1
M299 362 722 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=19120 $D=1
M300 359 355 361 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=14490 $D=1
M301 360 356 362 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=19120 $D=1
M302 361 57 229 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=14490 $D=1
M303 362 57 230 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=19120 $D=1
M304 233 58 361 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=14490 $D=1
M305 234 58 362 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=19120 $D=1
M306 363 58 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=14490 $D=1
M307 364 58 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=19120 $D=1
M308 6 59 365 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=14490 $D=1
M309 6 59 366 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=19120 $D=1
M310 367 60 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=14490 $D=1
M311 368 60 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=19120 $D=1
M312 369 59 219 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=14490 $D=1
M313 370 59 220 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=19120 $D=1
M314 6 369 723 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=14490 $D=1
M315 6 370 724 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=19120 $D=1
M316 371 723 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=14490 $D=1
M317 372 724 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=19120 $D=1
M318 369 365 371 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=14490 $D=1
M319 370 366 372 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=19120 $D=1
M320 371 60 229 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=14490 $D=1
M321 372 60 230 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=19120 $D=1
M322 233 61 371 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=14490 $D=1
M323 234 61 372 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=19120 $D=1
M324 373 61 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=14490 $D=1
M325 374 61 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=19120 $D=1
M326 6 62 375 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=14490 $D=1
M327 6 62 376 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=19120 $D=1
M328 377 63 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=14490 $D=1
M329 378 63 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=19120 $D=1
M330 379 62 219 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=14490 $D=1
M331 380 62 220 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=19120 $D=1
M332 6 379 725 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=14490 $D=1
M333 6 380 726 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=19120 $D=1
M334 381 725 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=14490 $D=1
M335 382 726 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=19120 $D=1
M336 379 375 381 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=14490 $D=1
M337 380 376 382 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=19120 $D=1
M338 381 63 229 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=14490 $D=1
M339 382 63 230 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=19120 $D=1
M340 233 64 381 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=14490 $D=1
M341 234 64 382 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=19120 $D=1
M342 383 64 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=14490 $D=1
M343 384 64 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=19120 $D=1
M344 6 65 385 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=14490 $D=1
M345 6 65 386 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=19120 $D=1
M346 387 66 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=14490 $D=1
M347 388 66 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=19120 $D=1
M348 389 65 219 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=14490 $D=1
M349 390 65 220 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=19120 $D=1
M350 6 389 727 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=14490 $D=1
M351 6 390 728 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=19120 $D=1
M352 391 727 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=14490 $D=1
M353 392 728 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=19120 $D=1
M354 389 385 391 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=14490 $D=1
M355 390 386 392 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=19120 $D=1
M356 391 66 229 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=14490 $D=1
M357 392 66 230 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=19120 $D=1
M358 233 67 391 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=14490 $D=1
M359 234 67 392 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=19120 $D=1
M360 393 67 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=14490 $D=1
M361 394 67 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=19120 $D=1
M362 6 68 395 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=14490 $D=1
M363 6 68 396 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=19120 $D=1
M364 397 69 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=14490 $D=1
M365 398 69 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=19120 $D=1
M366 399 68 219 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=14490 $D=1
M367 400 68 220 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=19120 $D=1
M368 6 399 729 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=14490 $D=1
M369 6 400 730 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=19120 $D=1
M370 401 729 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=14490 $D=1
M371 402 730 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=19120 $D=1
M372 399 395 401 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=14490 $D=1
M373 400 396 402 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=19120 $D=1
M374 401 69 229 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=14490 $D=1
M375 402 69 230 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=19120 $D=1
M376 233 70 401 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=14490 $D=1
M377 234 70 402 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=19120 $D=1
M378 403 70 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=14490 $D=1
M379 404 70 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=19120 $D=1
M380 6 71 405 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=14490 $D=1
M381 6 71 406 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=19120 $D=1
M382 407 72 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=14490 $D=1
M383 408 72 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=19120 $D=1
M384 409 71 219 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=14490 $D=1
M385 410 71 220 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=19120 $D=1
M386 6 409 731 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=14490 $D=1
M387 6 410 732 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=19120 $D=1
M388 411 731 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=14490 $D=1
M389 412 732 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=19120 $D=1
M390 409 405 411 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=14490 $D=1
M391 410 406 412 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=19120 $D=1
M392 411 72 229 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=14490 $D=1
M393 412 72 230 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=19120 $D=1
M394 233 73 411 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=14490 $D=1
M395 234 73 412 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=19120 $D=1
M396 413 73 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=14490 $D=1
M397 414 73 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=19120 $D=1
M398 6 74 415 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=14490 $D=1
M399 6 74 416 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=19120 $D=1
M400 417 75 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=14490 $D=1
M401 418 75 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=19120 $D=1
M402 419 74 219 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=14490 $D=1
M403 420 74 220 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=19120 $D=1
M404 6 419 733 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=14490 $D=1
M405 6 420 734 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=19120 $D=1
M406 421 733 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=14490 $D=1
M407 422 734 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=19120 $D=1
M408 419 415 421 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=14490 $D=1
M409 420 416 422 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=19120 $D=1
M410 421 75 229 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=14490 $D=1
M411 422 75 230 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=19120 $D=1
M412 233 76 421 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=14490 $D=1
M413 234 76 422 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=19120 $D=1
M414 423 76 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=14490 $D=1
M415 424 76 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=19120 $D=1
M416 6 77 425 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=14490 $D=1
M417 6 77 426 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=19120 $D=1
M418 427 78 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=14490 $D=1
M419 428 78 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=19120 $D=1
M420 429 77 219 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=14490 $D=1
M421 430 77 220 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=19120 $D=1
M422 6 429 735 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=14490 $D=1
M423 6 430 736 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=19120 $D=1
M424 431 735 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=14490 $D=1
M425 432 736 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=19120 $D=1
M426 429 425 431 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=14490 $D=1
M427 430 426 432 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=19120 $D=1
M428 431 78 229 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=14490 $D=1
M429 432 78 230 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=19120 $D=1
M430 233 79 431 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=14490 $D=1
M431 234 79 432 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=19120 $D=1
M432 433 79 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=14490 $D=1
M433 434 79 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=19120 $D=1
M434 6 80 435 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=14490 $D=1
M435 6 80 436 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=19120 $D=1
M436 437 81 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=14490 $D=1
M437 438 81 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=19120 $D=1
M438 439 80 219 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=14490 $D=1
M439 440 80 220 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=19120 $D=1
M440 6 439 737 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=14490 $D=1
M441 6 440 738 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=19120 $D=1
M442 441 737 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=14490 $D=1
M443 442 738 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=19120 $D=1
M444 439 435 441 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=14490 $D=1
M445 440 436 442 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=19120 $D=1
M446 441 81 229 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=14490 $D=1
M447 442 81 230 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=19120 $D=1
M448 233 82 441 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=14490 $D=1
M449 234 82 442 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=19120 $D=1
M450 443 82 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=14490 $D=1
M451 444 82 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=19120 $D=1
M452 6 83 445 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=14490 $D=1
M453 6 83 446 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=19120 $D=1
M454 447 84 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=14490 $D=1
M455 448 84 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=19120 $D=1
M456 449 83 219 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=14490 $D=1
M457 450 83 220 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=19120 $D=1
M458 6 449 739 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=14490 $D=1
M459 6 450 740 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=19120 $D=1
M460 451 739 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=14490 $D=1
M461 452 740 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=19120 $D=1
M462 449 445 451 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=14490 $D=1
M463 450 446 452 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=19120 $D=1
M464 451 84 229 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=14490 $D=1
M465 452 84 230 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=19120 $D=1
M466 233 85 451 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=14490 $D=1
M467 234 85 452 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=19120 $D=1
M468 453 85 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=14490 $D=1
M469 454 85 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=19120 $D=1
M470 6 86 455 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=14490 $D=1
M471 6 86 456 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=19120 $D=1
M472 457 87 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=14490 $D=1
M473 458 87 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=19120 $D=1
M474 459 86 219 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=14490 $D=1
M475 460 86 220 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=19120 $D=1
M476 6 459 741 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=14490 $D=1
M477 6 460 742 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=19120 $D=1
M478 461 741 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=14490 $D=1
M479 462 742 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=19120 $D=1
M480 459 455 461 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=14490 $D=1
M481 460 456 462 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=19120 $D=1
M482 461 87 229 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=14490 $D=1
M483 462 87 230 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=19120 $D=1
M484 233 88 461 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=14490 $D=1
M485 234 88 462 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=19120 $D=1
M486 463 88 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=14490 $D=1
M487 464 88 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=19120 $D=1
M488 6 89 465 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=14490 $D=1
M489 6 89 466 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=19120 $D=1
M490 467 90 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=14490 $D=1
M491 468 90 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=19120 $D=1
M492 469 89 219 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=14490 $D=1
M493 470 89 220 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=19120 $D=1
M494 6 469 743 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=14490 $D=1
M495 6 470 744 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=19120 $D=1
M496 471 743 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=14490 $D=1
M497 472 744 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=19120 $D=1
M498 469 465 471 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=14490 $D=1
M499 470 466 472 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=19120 $D=1
M500 471 90 229 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=14490 $D=1
M501 472 90 230 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=19120 $D=1
M502 233 91 471 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=14490 $D=1
M503 234 91 472 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=19120 $D=1
M504 473 91 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=14490 $D=1
M505 474 91 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=19120 $D=1
M506 6 92 475 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=14490 $D=1
M507 6 92 476 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=19120 $D=1
M508 477 93 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=14490 $D=1
M509 478 93 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=19120 $D=1
M510 479 92 219 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=14490 $D=1
M511 480 92 220 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=19120 $D=1
M512 6 479 745 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=14490 $D=1
M513 6 480 746 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=19120 $D=1
M514 481 745 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=14490 $D=1
M515 482 746 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=19120 $D=1
M516 479 475 481 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=14490 $D=1
M517 480 476 482 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=19120 $D=1
M518 481 93 229 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=14490 $D=1
M519 482 93 230 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=19120 $D=1
M520 233 94 481 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=14490 $D=1
M521 234 94 482 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=19120 $D=1
M522 483 94 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=14490 $D=1
M523 484 94 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=19120 $D=1
M524 6 95 485 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=14490 $D=1
M525 6 95 486 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=19120 $D=1
M526 487 96 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=14490 $D=1
M527 488 96 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=19120 $D=1
M528 489 95 219 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=14490 $D=1
M529 490 95 220 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=19120 $D=1
M530 6 489 747 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=14490 $D=1
M531 6 490 748 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=19120 $D=1
M532 491 747 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=14490 $D=1
M533 492 748 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=19120 $D=1
M534 489 485 491 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=14490 $D=1
M535 490 486 492 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=19120 $D=1
M536 491 96 229 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=14490 $D=1
M537 492 96 230 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=19120 $D=1
M538 233 97 491 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=14490 $D=1
M539 234 97 492 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=19120 $D=1
M540 493 97 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=14490 $D=1
M541 494 97 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=19120 $D=1
M542 6 98 495 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=14490 $D=1
M543 6 98 496 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=19120 $D=1
M544 497 99 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=14490 $D=1
M545 498 99 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=19120 $D=1
M546 499 98 219 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=14490 $D=1
M547 500 98 220 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=19120 $D=1
M548 6 499 749 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=14490 $D=1
M549 6 500 750 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=19120 $D=1
M550 501 749 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=14490 $D=1
M551 502 750 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=19120 $D=1
M552 499 495 501 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=14490 $D=1
M553 500 496 502 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=19120 $D=1
M554 501 99 229 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=14490 $D=1
M555 502 99 230 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=19120 $D=1
M556 233 100 501 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=14490 $D=1
M557 234 100 502 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=19120 $D=1
M558 503 100 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=14490 $D=1
M559 504 100 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=19120 $D=1
M560 6 101 505 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=14490 $D=1
M561 6 101 506 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=19120 $D=1
M562 507 102 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=14490 $D=1
M563 508 102 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=19120 $D=1
M564 509 101 219 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=14490 $D=1
M565 510 101 220 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=19120 $D=1
M566 6 509 751 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=14490 $D=1
M567 6 510 752 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=19120 $D=1
M568 511 751 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=14490 $D=1
M569 512 752 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=19120 $D=1
M570 509 505 511 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=14490 $D=1
M571 510 506 512 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=19120 $D=1
M572 511 102 229 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=14490 $D=1
M573 512 102 230 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=19120 $D=1
M574 233 103 511 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=14490 $D=1
M575 234 103 512 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=19120 $D=1
M576 513 103 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=14490 $D=1
M577 514 103 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=19120 $D=1
M578 6 104 515 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=14490 $D=1
M579 6 104 516 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=19120 $D=1
M580 517 105 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=14490 $D=1
M581 518 105 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=19120 $D=1
M582 519 104 219 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=14490 $D=1
M583 520 104 220 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=19120 $D=1
M584 6 519 753 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=14490 $D=1
M585 6 520 754 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=19120 $D=1
M586 521 753 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=14490 $D=1
M587 522 754 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=19120 $D=1
M588 519 515 521 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=14490 $D=1
M589 520 516 522 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=19120 $D=1
M590 521 105 229 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=14490 $D=1
M591 522 105 230 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=19120 $D=1
M592 233 107 521 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=14490 $D=1
M593 234 107 522 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=19120 $D=1
M594 523 107 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=14490 $D=1
M595 524 107 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=19120 $D=1
M596 6 109 525 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=14490 $D=1
M597 6 109 526 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=19120 $D=1
M598 527 110 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=14490 $D=1
M599 528 110 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=19120 $D=1
M600 529 109 219 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=14490 $D=1
M601 530 109 220 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=19120 $D=1
M602 6 529 755 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=14490 $D=1
M603 6 530 756 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=19120 $D=1
M604 531 755 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=14490 $D=1
M605 532 756 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=19120 $D=1
M606 529 525 531 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=14490 $D=1
M607 530 526 532 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=19120 $D=1
M608 531 110 229 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=14490 $D=1
M609 532 110 230 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=19120 $D=1
M610 233 113 531 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=14490 $D=1
M611 234 113 532 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=19120 $D=1
M612 533 113 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=14490 $D=1
M613 534 113 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=19120 $D=1
M614 6 114 535 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=14490 $D=1
M615 6 114 536 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=19120 $D=1
M616 537 115 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=14490 $D=1
M617 538 115 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=19120 $D=1
M618 6 115 229 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=14490 $D=1
M619 6 115 230 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=19120 $D=1
M620 233 114 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=14490 $D=1
M621 234 114 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=19120 $D=1
M622 6 541 539 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=14490 $D=1
M623 6 542 540 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=19120 $D=1
M624 541 116 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=14490 $D=1
M625 542 116 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=19120 $D=1
M626 757 229 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=14490 $D=1
M627 758 230 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=19120 $D=1
M628 543 539 757 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=14490 $D=1
M629 544 540 758 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=19120 $D=1
M630 6 543 545 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=14490 $D=1
M631 6 544 546 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=19120 $D=1
M632 759 545 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=14490 $D=1
M633 760 546 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=19120 $D=1
M634 543 541 759 6 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=14490 $D=1
M635 544 542 760 6 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=19120 $D=1
M636 6 549 547 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=14490 $D=1
M637 6 550 548 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=19120 $D=1
M638 549 116 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=14490 $D=1
M639 550 116 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=19120 $D=1
M640 761 233 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=14490 $D=1
M641 762 234 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=19120 $D=1
M642 551 547 761 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=14490 $D=1
M643 552 548 762 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=19120 $D=1
M644 6 551 117 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=14490 $D=1
M645 6 552 118 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=19120 $D=1
M646 763 117 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=14490 $D=1
M647 764 118 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=19120 $D=1
M648 551 549 763 6 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=14490 $D=1
M649 552 550 764 6 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=19120 $D=1
M650 553 119 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=14490 $D=1
M651 554 119 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=19120 $D=1
M652 555 553 545 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=14490 $D=1
M653 556 554 546 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=19120 $D=1
M654 120 119 555 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=14490 $D=1
M655 121 119 556 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=19120 $D=1
M656 557 122 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=14490 $D=1
M657 558 122 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=19120 $D=1
M658 559 557 117 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=14490 $D=1
M659 560 558 118 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=19120 $D=1
M660 765 122 559 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=14490 $D=1
M661 766 122 560 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=19120 $D=1
M662 6 117 765 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=14490 $D=1
M663 6 118 766 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=19120 $D=1
M664 561 123 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=14490 $D=1
M665 562 123 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=19120 $D=1
M666 563 561 559 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=14490 $D=1
M667 564 562 560 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=19120 $D=1
M668 11 123 563 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=14490 $D=1
M669 12 123 564 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=19120 $D=1
M670 566 565 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=14490 $D=1
M671 567 124 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=19120 $D=1
M672 6 570 568 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=14490 $D=1
M673 6 571 569 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=19120 $D=1
M674 572 555 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=14490 $D=1
M675 573 556 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=19120 $D=1
M676 570 572 565 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=14490 $D=1
M677 571 573 124 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=19120 $D=1
M678 566 555 570 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=14490 $D=1
M679 567 556 571 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=19120 $D=1
M680 574 568 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=14490 $D=1
M681 575 569 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=19120 $D=1
M682 125 574 563 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=14490 $D=1
M683 565 575 564 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=19120 $D=1
M684 555 568 125 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=14490 $D=1
M685 556 569 565 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=19120 $D=1
M686 576 125 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=14490 $D=1
M687 577 565 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=19120 $D=1
M688 578 568 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=14490 $D=1
M689 579 569 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=19120 $D=1
M690 580 578 576 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=14490 $D=1
M691 581 579 577 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=19120 $D=1
M692 563 568 580 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=14490 $D=1
M693 564 569 581 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=19120 $D=1
M694 582 555 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=14490 $D=1
M695 583 556 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=19120 $D=1
M696 6 563 582 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=14490 $D=1
M697 6 564 583 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=19120 $D=1
M698 584 580 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=14490 $D=1
M699 585 581 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=19120 $D=1
M700 785 555 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=14490 $D=1
M701 786 556 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=19120 $D=1
M702 586 563 785 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=14490 $D=1
M703 587 564 786 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=19120 $D=1
M704 787 555 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=14490 $D=1
M705 788 556 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=19120 $D=1
M706 588 563 787 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=14490 $D=1
M707 589 564 788 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=19120 $D=1
M708 592 555 590 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=14490 $D=1
M709 593 556 591 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=19120 $D=1
M710 590 563 592 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=14490 $D=1
M711 591 564 593 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=19120 $D=1
M712 6 588 590 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=14490 $D=1
M713 6 589 591 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=19120 $D=1
M714 594 128 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=14490 $D=1
M715 595 128 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=19120 $D=1
M716 596 594 582 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=14490 $D=1
M717 597 595 583 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=19120 $D=1
M718 586 128 596 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=14490 $D=1
M719 587 128 597 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=19120 $D=1
M720 598 594 584 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=14490 $D=1
M721 599 595 585 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=19120 $D=1
M722 592 128 598 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=14490 $D=1
M723 593 128 599 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=19120 $D=1
M724 600 129 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=14490 $D=1
M725 601 129 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=19120 $D=1
M726 602 600 598 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=14490 $D=1
M727 603 601 599 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=19120 $D=1
M728 596 129 602 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=14490 $D=1
M729 597 129 603 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=19120 $D=1
M730 13 602 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=14490 $D=1
M731 14 603 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=19120 $D=1
M732 604 130 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=14490 $D=1
M733 605 130 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=19120 $D=1
M734 606 604 131 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=14490 $D=1
M735 607 605 132 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=19120 $D=1
M736 133 130 606 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=14490 $D=1
M737 134 130 607 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=19120 $D=1
M738 608 130 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=14490 $D=1
M739 609 130 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=19120 $D=1
M740 610 608 135 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=14490 $D=1
M741 611 609 136 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=19120 $D=1
M742 137 130 610 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=14490 $D=1
M743 138 130 611 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=19120 $D=1
M744 612 130 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=14490 $D=1
M745 613 130 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=19120 $D=1
M746 614 612 126 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=14490 $D=1
M747 615 613 127 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=19120 $D=1
M748 139 130 614 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=14490 $D=1
M749 140 130 615 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=19120 $D=1
M750 616 130 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=14490 $D=1
M751 617 130 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=19120 $D=1
M752 618 616 142 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=14490 $D=1
M753 619 617 143 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=19120 $D=1
M754 139 130 618 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=14490 $D=1
M755 139 130 619 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=19120 $D=1
M756 620 130 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=14490 $D=1
M757 621 130 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=19120 $D=1
M758 622 620 144 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=14490 $D=1
M759 623 621 145 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=19120 $D=1
M760 139 130 622 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=14490 $D=1
M761 139 130 623 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=19120 $D=1
M762 6 555 767 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=14490 $D=1
M763 6 556 768 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=19120 $D=1
M764 134 767 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=14490 $D=1
M765 131 768 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=19120 $D=1
M766 624 146 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=14490 $D=1
M767 625 146 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=19120 $D=1
M768 147 624 134 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=14490 $D=1
M769 148 625 131 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=19120 $D=1
M770 606 146 147 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=14490 $D=1
M771 607 146 148 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=19120 $D=1
M772 626 149 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=14490 $D=1
M773 627 149 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=19120 $D=1
M774 150 626 147 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=14490 $D=1
M775 106 627 148 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=19120 $D=1
M776 610 149 150 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=14490 $D=1
M777 611 149 106 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=19120 $D=1
M778 628 151 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=14490 $D=1
M779 629 151 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=19120 $D=1
M780 152 628 150 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=14490 $D=1
M781 111 629 106 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=19120 $D=1
M782 614 151 152 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=14490 $D=1
M783 615 151 111 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=19120 $D=1
M784 630 153 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=14490 $D=1
M785 631 153 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=19120 $D=1
M786 154 630 152 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=14490 $D=1
M787 155 631 111 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=19120 $D=1
M788 618 153 154 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=14490 $D=1
M789 619 153 155 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=19120 $D=1
M790 632 156 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=14490 $D=1
M791 633 156 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=19120 $D=1
M792 205 632 154 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=14490 $D=1
M793 206 633 155 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=19120 $D=1
M794 622 156 205 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=14490 $D=1
M795 623 156 206 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=19120 $D=1
M796 634 157 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=14490 $D=1
M797 635 157 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=19120 $D=1
M798 636 634 117 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=14490 $D=1
M799 637 635 118 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=19120 $D=1
M800 11 157 636 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=14490 $D=1
M801 12 157 637 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=19120 $D=1
M802 789 545 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=14490 $D=1
M803 790 546 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=19120 $D=1
M804 638 636 789 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=14490 $D=1
M805 639 637 790 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=19120 $D=1
M806 642 545 640 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=14490 $D=1
M807 643 546 641 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=19120 $D=1
M808 640 636 642 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=14490 $D=1
M809 641 637 643 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=19120 $D=1
M810 6 638 640 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=14490 $D=1
M811 6 639 641 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=19120 $D=1
M812 791 158 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=14490 $D=1
M813 792 644 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=19120 $D=1
M814 769 642 791 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=14490 $D=1
M815 770 643 792 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=19120 $D=1
M816 644 769 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=14490 $D=1
M817 159 770 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=19120 $D=1
M818 645 545 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=14490 $D=1
M819 646 546 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=19120 $D=1
M820 6 647 645 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=14490 $D=1
M821 6 648 646 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=19120 $D=1
M822 647 636 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=14490 $D=1
M823 648 637 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=19120 $D=1
M824 793 645 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=14490 $D=1
M825 794 646 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=19120 $D=1
M826 649 158 793 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=14490 $D=1
M827 650 644 794 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=19120 $D=1
M828 652 160 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=14490 $D=1
M829 653 651 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=19120 $D=1
M830 795 649 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=14490 $D=1
M831 796 650 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=19120 $D=1
M832 651 652 795 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=14490 $D=1
M833 161 653 796 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=19120 $D=1
M834 655 654 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=14490 $D=1
M835 656 162 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=19120 $D=1
M836 6 659 657 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=14490 $D=1
M837 6 660 658 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=19120 $D=1
M838 661 120 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=14490 $D=1
M839 662 121 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=19120 $D=1
M840 659 661 654 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=14490 $D=1
M841 660 662 162 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=19120 $D=1
M842 655 120 659 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=14490 $D=1
M843 656 121 660 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=19120 $D=1
M844 663 657 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=14490 $D=1
M845 664 658 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=19120 $D=1
M846 163 663 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=14490 $D=1
M847 654 664 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=19120 $D=1
M848 120 657 163 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=14490 $D=1
M849 121 658 654 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=19120 $D=1
M850 665 163 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=14490 $D=1
M851 666 654 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=19120 $D=1
M852 667 657 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=14490 $D=1
M853 668 658 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=19120 $D=1
M854 207 667 665 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=14490 $D=1
M855 208 668 666 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=19120 $D=1
M856 6 657 207 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=14490 $D=1
M857 6 658 208 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=19120 $D=1
M858 669 164 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=14490 $D=1
M859 670 164 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=19120 $D=1
M860 671 669 207 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=14490 $D=1
M861 672 670 208 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=19120 $D=1
M862 13 164 671 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=14490 $D=1
M863 14 164 672 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=19120 $D=1
M864 673 165 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=14490 $D=1
M865 674 165 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=19120 $D=1
M866 675 673 671 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=14490 $D=1
M867 676 674 672 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=19120 $D=1
M868 6 165 675 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=14490 $D=1
M869 6 165 676 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=19120 $D=1
M870 677 116 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=14490 $D=1
M871 678 116 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=19120 $D=1
M872 6 677 679 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=14490 $D=1
M873 6 678 680 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=19120 $D=1
M874 681 116 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=14490 $D=1
M875 682 116 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=19120 $D=1
M876 683 677 675 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=14490 $D=1
M877 684 678 676 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=19120 $D=1
M878 6 683 771 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=14490 $D=1
M879 6 684 772 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=19120 $D=1
M880 685 771 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=14490 $D=1
M881 686 772 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=19120 $D=1
M882 683 679 685 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=14490 $D=1
M883 684 680 686 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=19120 $D=1
M884 687 116 685 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=14490 $D=1
M885 688 116 686 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=19120 $D=1
M886 6 691 689 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=14490 $D=1
M887 6 692 690 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=19120 $D=1
M888 691 116 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=14490 $D=1
M889 692 116 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=19120 $D=1
M890 773 687 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=14490 $D=1
M891 774 688 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=19120 $D=1
M892 693 689 773 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=14490 $D=1
M893 694 690 774 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=19120 $D=1
M894 6 693 120 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=14490 $D=1
M895 6 694 121 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=19120 $D=1
M896 775 120 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=14490 $D=1
M897 776 121 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=19120 $D=1
M898 693 691 775 6 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=14490 $D=1
M899 694 692 776 6 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=19120 $D=1
M900 181 1 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=15740 $D=0
M901 182 1 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=20370 $D=0
M902 183 1 2 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=15740 $D=0
M903 184 1 3 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=20370 $D=0
M904 6 181 183 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=15740 $D=0
M905 6 182 184 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=20370 $D=0
M906 185 1 4 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=15740 $D=0
M907 186 1 4 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=20370 $D=0
M908 5 181 185 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=15740 $D=0
M909 5 182 186 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=20370 $D=0
M910 187 1 6 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=15740 $D=0
M911 188 1 6 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=20370 $D=0
M912 6 181 187 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=15740 $D=0
M913 6 182 188 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=20370 $D=0
M914 191 7 187 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=15740 $D=0
M915 192 7 188 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=20370 $D=0
M916 189 7 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=15740 $D=0
M917 190 7 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=20370 $D=0
M918 193 7 185 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=15740 $D=0
M919 194 7 186 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=20370 $D=0
M920 183 189 193 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=15740 $D=0
M921 184 190 194 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=20370 $D=0
M922 195 8 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=15740 $D=0
M923 196 8 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=20370 $D=0
M924 197 8 193 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=15740 $D=0
M925 198 8 194 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=20370 $D=0
M926 191 195 197 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=15740 $D=0
M927 192 196 198 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=20370 $D=0
M928 199 10 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=15740 $D=0
M929 200 10 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=20370 $D=0
M930 201 10 6 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=15740 $D=0
M931 202 10 6 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=20370 $D=0
M932 11 199 201 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=15740 $D=0
M933 12 200 202 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=20370 $D=0
M934 203 10 13 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=15740 $D=0
M935 204 10 14 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=20370 $D=0
M936 205 199 203 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=15740 $D=0
M937 206 200 204 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=20370 $D=0
M938 209 10 207 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=15740 $D=0
M939 210 10 208 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=20370 $D=0
M940 197 199 209 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=15740 $D=0
M941 198 200 210 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=20370 $D=0
M942 213 15 209 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=15740 $D=0
M943 214 15 210 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=20370 $D=0
M944 211 15 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=15740 $D=0
M945 212 15 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=20370 $D=0
M946 215 15 203 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=15740 $D=0
M947 216 15 204 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=20370 $D=0
M948 201 211 215 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=15740 $D=0
M949 202 212 216 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=20370 $D=0
M950 217 16 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=15740 $D=0
M951 218 16 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=20370 $D=0
M952 219 16 215 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=15740 $D=0
M953 220 16 216 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=20370 $D=0
M954 213 217 219 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=15740 $D=0
M955 214 218 220 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=20370 $D=0
M956 9 17 221 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=15740 $D=0
M957 9 17 222 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=20370 $D=0
M958 223 18 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=15740 $D=0
M959 224 18 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=20370 $D=0
M960 225 221 219 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=15740 $D=0
M961 226 222 220 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=20370 $D=0
M962 9 225 695 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=15740 $D=0
M963 9 226 696 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=20370 $D=0
M964 227 695 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=15740 $D=0
M965 228 696 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=20370 $D=0
M966 225 17 227 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=15740 $D=0
M967 226 17 228 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=20370 $D=0
M968 227 223 229 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=15740 $D=0
M969 228 224 230 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=20370 $D=0
M970 233 231 227 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=15740 $D=0
M971 234 232 228 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=20370 $D=0
M972 231 19 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=15740 $D=0
M973 232 19 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=20370 $D=0
M974 9 20 235 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=15740 $D=0
M975 9 20 236 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=20370 $D=0
M976 237 21 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=15740 $D=0
M977 238 21 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=20370 $D=0
M978 239 235 219 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=15740 $D=0
M979 240 236 220 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=20370 $D=0
M980 9 239 697 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=15740 $D=0
M981 9 240 698 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=20370 $D=0
M982 241 697 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=15740 $D=0
M983 242 698 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=20370 $D=0
M984 239 20 241 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=15740 $D=0
M985 240 20 242 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=20370 $D=0
M986 241 237 229 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=15740 $D=0
M987 242 238 230 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=20370 $D=0
M988 233 243 241 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=15740 $D=0
M989 234 244 242 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=20370 $D=0
M990 243 22 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=15740 $D=0
M991 244 22 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=20370 $D=0
M992 9 23 245 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=15740 $D=0
M993 9 23 246 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=20370 $D=0
M994 247 24 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=15740 $D=0
M995 248 24 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=20370 $D=0
M996 249 245 219 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=15740 $D=0
M997 250 246 220 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=20370 $D=0
M998 9 249 699 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=15740 $D=0
M999 9 250 700 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=20370 $D=0
M1000 251 699 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=15740 $D=0
M1001 252 700 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=20370 $D=0
M1002 249 23 251 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=15740 $D=0
M1003 250 23 252 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=20370 $D=0
M1004 251 247 229 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=15740 $D=0
M1005 252 248 230 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=20370 $D=0
M1006 233 253 251 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=15740 $D=0
M1007 234 254 252 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=20370 $D=0
M1008 253 25 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=15740 $D=0
M1009 254 25 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=20370 $D=0
M1010 9 26 255 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=15740 $D=0
M1011 9 26 256 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=20370 $D=0
M1012 257 27 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=15740 $D=0
M1013 258 27 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=20370 $D=0
M1014 259 255 219 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=15740 $D=0
M1015 260 256 220 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=20370 $D=0
M1016 9 259 701 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=15740 $D=0
M1017 9 260 702 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=20370 $D=0
M1018 261 701 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=15740 $D=0
M1019 262 702 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=20370 $D=0
M1020 259 26 261 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=15740 $D=0
M1021 260 26 262 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=20370 $D=0
M1022 261 257 229 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=15740 $D=0
M1023 262 258 230 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=20370 $D=0
M1024 233 263 261 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=15740 $D=0
M1025 234 264 262 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=20370 $D=0
M1026 263 28 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=15740 $D=0
M1027 264 28 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=20370 $D=0
M1028 9 29 265 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=15740 $D=0
M1029 9 29 266 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=20370 $D=0
M1030 267 30 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=15740 $D=0
M1031 268 30 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=20370 $D=0
M1032 269 265 219 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=15740 $D=0
M1033 270 266 220 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=20370 $D=0
M1034 9 269 703 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=15740 $D=0
M1035 9 270 704 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=20370 $D=0
M1036 271 703 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=15740 $D=0
M1037 272 704 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=20370 $D=0
M1038 269 29 271 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=15740 $D=0
M1039 270 29 272 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=20370 $D=0
M1040 271 267 229 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=15740 $D=0
M1041 272 268 230 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=20370 $D=0
M1042 233 273 271 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=15740 $D=0
M1043 234 274 272 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=20370 $D=0
M1044 273 31 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=15740 $D=0
M1045 274 31 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=20370 $D=0
M1046 9 32 275 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=15740 $D=0
M1047 9 32 276 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=20370 $D=0
M1048 277 33 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=15740 $D=0
M1049 278 33 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=20370 $D=0
M1050 279 275 219 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=15740 $D=0
M1051 280 276 220 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=20370 $D=0
M1052 9 279 705 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=15740 $D=0
M1053 9 280 706 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=20370 $D=0
M1054 281 705 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=15740 $D=0
M1055 282 706 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=20370 $D=0
M1056 279 32 281 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=15740 $D=0
M1057 280 32 282 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=20370 $D=0
M1058 281 277 229 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=15740 $D=0
M1059 282 278 230 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=20370 $D=0
M1060 233 283 281 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=15740 $D=0
M1061 234 284 282 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=20370 $D=0
M1062 283 34 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=15740 $D=0
M1063 284 34 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=20370 $D=0
M1064 9 35 285 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=15740 $D=0
M1065 9 35 286 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=20370 $D=0
M1066 287 36 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=15740 $D=0
M1067 288 36 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=20370 $D=0
M1068 289 285 219 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=15740 $D=0
M1069 290 286 220 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=20370 $D=0
M1070 9 289 707 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=15740 $D=0
M1071 9 290 708 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=20370 $D=0
M1072 291 707 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=15740 $D=0
M1073 292 708 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=20370 $D=0
M1074 289 35 291 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=15740 $D=0
M1075 290 35 292 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=20370 $D=0
M1076 291 287 229 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=15740 $D=0
M1077 292 288 230 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=20370 $D=0
M1078 233 293 291 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=15740 $D=0
M1079 234 294 292 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=20370 $D=0
M1080 293 37 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=15740 $D=0
M1081 294 37 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=20370 $D=0
M1082 9 38 295 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=15740 $D=0
M1083 9 38 296 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=20370 $D=0
M1084 297 39 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=15740 $D=0
M1085 298 39 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=20370 $D=0
M1086 299 295 219 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=15740 $D=0
M1087 300 296 220 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=20370 $D=0
M1088 9 299 709 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=15740 $D=0
M1089 9 300 710 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=20370 $D=0
M1090 301 709 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=15740 $D=0
M1091 302 710 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=20370 $D=0
M1092 299 38 301 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=15740 $D=0
M1093 300 38 302 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=20370 $D=0
M1094 301 297 229 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=15740 $D=0
M1095 302 298 230 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=20370 $D=0
M1096 233 303 301 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=15740 $D=0
M1097 234 304 302 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=20370 $D=0
M1098 303 40 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=15740 $D=0
M1099 304 40 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=20370 $D=0
M1100 9 41 305 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=15740 $D=0
M1101 9 41 306 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=20370 $D=0
M1102 307 42 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=15740 $D=0
M1103 308 42 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=20370 $D=0
M1104 309 305 219 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=15740 $D=0
M1105 310 306 220 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=20370 $D=0
M1106 9 309 711 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=15740 $D=0
M1107 9 310 712 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=20370 $D=0
M1108 311 711 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=15740 $D=0
M1109 312 712 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=20370 $D=0
M1110 309 41 311 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=15740 $D=0
M1111 310 41 312 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=20370 $D=0
M1112 311 307 229 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=15740 $D=0
M1113 312 308 230 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=20370 $D=0
M1114 233 313 311 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=15740 $D=0
M1115 234 314 312 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=20370 $D=0
M1116 313 43 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=15740 $D=0
M1117 314 43 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=20370 $D=0
M1118 9 44 315 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=15740 $D=0
M1119 9 44 316 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=20370 $D=0
M1120 317 45 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=15740 $D=0
M1121 318 45 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=20370 $D=0
M1122 319 315 219 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=15740 $D=0
M1123 320 316 220 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=20370 $D=0
M1124 9 319 713 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=15740 $D=0
M1125 9 320 714 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=20370 $D=0
M1126 321 713 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=15740 $D=0
M1127 322 714 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=20370 $D=0
M1128 319 44 321 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=15740 $D=0
M1129 320 44 322 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=20370 $D=0
M1130 321 317 229 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=15740 $D=0
M1131 322 318 230 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=20370 $D=0
M1132 233 323 321 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=15740 $D=0
M1133 234 324 322 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=20370 $D=0
M1134 323 46 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=15740 $D=0
M1135 324 46 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=20370 $D=0
M1136 9 47 325 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=15740 $D=0
M1137 9 47 326 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=20370 $D=0
M1138 327 48 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=15740 $D=0
M1139 328 48 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=20370 $D=0
M1140 329 325 219 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=15740 $D=0
M1141 330 326 220 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=20370 $D=0
M1142 9 329 715 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=15740 $D=0
M1143 9 330 716 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=20370 $D=0
M1144 331 715 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=15740 $D=0
M1145 332 716 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=20370 $D=0
M1146 329 47 331 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=15740 $D=0
M1147 330 47 332 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=20370 $D=0
M1148 331 327 229 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=15740 $D=0
M1149 332 328 230 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=20370 $D=0
M1150 233 333 331 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=15740 $D=0
M1151 234 334 332 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=20370 $D=0
M1152 333 49 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=15740 $D=0
M1153 334 49 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=20370 $D=0
M1154 9 50 335 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=15740 $D=0
M1155 9 50 336 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=20370 $D=0
M1156 337 51 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=15740 $D=0
M1157 338 51 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=20370 $D=0
M1158 339 335 219 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=15740 $D=0
M1159 340 336 220 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=20370 $D=0
M1160 9 339 717 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=15740 $D=0
M1161 9 340 718 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=20370 $D=0
M1162 341 717 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=15740 $D=0
M1163 342 718 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=20370 $D=0
M1164 339 50 341 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=15740 $D=0
M1165 340 50 342 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=20370 $D=0
M1166 341 337 229 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=15740 $D=0
M1167 342 338 230 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=20370 $D=0
M1168 233 343 341 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=15740 $D=0
M1169 234 344 342 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=20370 $D=0
M1170 343 52 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=15740 $D=0
M1171 344 52 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=20370 $D=0
M1172 9 53 345 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=15740 $D=0
M1173 9 53 346 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=20370 $D=0
M1174 347 54 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=15740 $D=0
M1175 348 54 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=20370 $D=0
M1176 349 345 219 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=15740 $D=0
M1177 350 346 220 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=20370 $D=0
M1178 9 349 719 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=15740 $D=0
M1179 9 350 720 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=20370 $D=0
M1180 351 719 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=15740 $D=0
M1181 352 720 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=20370 $D=0
M1182 349 53 351 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=15740 $D=0
M1183 350 53 352 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=20370 $D=0
M1184 351 347 229 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=15740 $D=0
M1185 352 348 230 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=20370 $D=0
M1186 233 353 351 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=15740 $D=0
M1187 234 354 352 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=20370 $D=0
M1188 353 55 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=15740 $D=0
M1189 354 55 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=20370 $D=0
M1190 9 56 355 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=15740 $D=0
M1191 9 56 356 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=20370 $D=0
M1192 357 57 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=15740 $D=0
M1193 358 57 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=20370 $D=0
M1194 359 355 219 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=15740 $D=0
M1195 360 356 220 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=20370 $D=0
M1196 9 359 721 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=15740 $D=0
M1197 9 360 722 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=20370 $D=0
M1198 361 721 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=15740 $D=0
M1199 362 722 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=20370 $D=0
M1200 359 56 361 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=15740 $D=0
M1201 360 56 362 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=20370 $D=0
M1202 361 357 229 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=15740 $D=0
M1203 362 358 230 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=20370 $D=0
M1204 233 363 361 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=15740 $D=0
M1205 234 364 362 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=20370 $D=0
M1206 363 58 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=15740 $D=0
M1207 364 58 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=20370 $D=0
M1208 9 59 365 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=15740 $D=0
M1209 9 59 366 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=20370 $D=0
M1210 367 60 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=15740 $D=0
M1211 368 60 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=20370 $D=0
M1212 369 365 219 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=15740 $D=0
M1213 370 366 220 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=20370 $D=0
M1214 9 369 723 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=15740 $D=0
M1215 9 370 724 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=20370 $D=0
M1216 371 723 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=15740 $D=0
M1217 372 724 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=20370 $D=0
M1218 369 59 371 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=15740 $D=0
M1219 370 59 372 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=20370 $D=0
M1220 371 367 229 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=15740 $D=0
M1221 372 368 230 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=20370 $D=0
M1222 233 373 371 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=15740 $D=0
M1223 234 374 372 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=20370 $D=0
M1224 373 61 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=15740 $D=0
M1225 374 61 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=20370 $D=0
M1226 9 62 375 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=15740 $D=0
M1227 9 62 376 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=20370 $D=0
M1228 377 63 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=15740 $D=0
M1229 378 63 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=20370 $D=0
M1230 379 375 219 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=15740 $D=0
M1231 380 376 220 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=20370 $D=0
M1232 9 379 725 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=15740 $D=0
M1233 9 380 726 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=20370 $D=0
M1234 381 725 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=15740 $D=0
M1235 382 726 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=20370 $D=0
M1236 379 62 381 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=15740 $D=0
M1237 380 62 382 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=20370 $D=0
M1238 381 377 229 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=15740 $D=0
M1239 382 378 230 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=20370 $D=0
M1240 233 383 381 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=15740 $D=0
M1241 234 384 382 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=20370 $D=0
M1242 383 64 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=15740 $D=0
M1243 384 64 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=20370 $D=0
M1244 9 65 385 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=15740 $D=0
M1245 9 65 386 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=20370 $D=0
M1246 387 66 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=15740 $D=0
M1247 388 66 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=20370 $D=0
M1248 389 385 219 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=15740 $D=0
M1249 390 386 220 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=20370 $D=0
M1250 9 389 727 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=15740 $D=0
M1251 9 390 728 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=20370 $D=0
M1252 391 727 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=15740 $D=0
M1253 392 728 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=20370 $D=0
M1254 389 65 391 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=15740 $D=0
M1255 390 65 392 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=20370 $D=0
M1256 391 387 229 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=15740 $D=0
M1257 392 388 230 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=20370 $D=0
M1258 233 393 391 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=15740 $D=0
M1259 234 394 392 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=20370 $D=0
M1260 393 67 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=15740 $D=0
M1261 394 67 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=20370 $D=0
M1262 9 68 395 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=15740 $D=0
M1263 9 68 396 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=20370 $D=0
M1264 397 69 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=15740 $D=0
M1265 398 69 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=20370 $D=0
M1266 399 395 219 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=15740 $D=0
M1267 400 396 220 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=20370 $D=0
M1268 9 399 729 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=15740 $D=0
M1269 9 400 730 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=20370 $D=0
M1270 401 729 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=15740 $D=0
M1271 402 730 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=20370 $D=0
M1272 399 68 401 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=15740 $D=0
M1273 400 68 402 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=20370 $D=0
M1274 401 397 229 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=15740 $D=0
M1275 402 398 230 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=20370 $D=0
M1276 233 403 401 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=15740 $D=0
M1277 234 404 402 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=20370 $D=0
M1278 403 70 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=15740 $D=0
M1279 404 70 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=20370 $D=0
M1280 9 71 405 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=15740 $D=0
M1281 9 71 406 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=20370 $D=0
M1282 407 72 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=15740 $D=0
M1283 408 72 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=20370 $D=0
M1284 409 405 219 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=15740 $D=0
M1285 410 406 220 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=20370 $D=0
M1286 9 409 731 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=15740 $D=0
M1287 9 410 732 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=20370 $D=0
M1288 411 731 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=15740 $D=0
M1289 412 732 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=20370 $D=0
M1290 409 71 411 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=15740 $D=0
M1291 410 71 412 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=20370 $D=0
M1292 411 407 229 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=15740 $D=0
M1293 412 408 230 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=20370 $D=0
M1294 233 413 411 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=15740 $D=0
M1295 234 414 412 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=20370 $D=0
M1296 413 73 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=15740 $D=0
M1297 414 73 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=20370 $D=0
M1298 9 74 415 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=15740 $D=0
M1299 9 74 416 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=20370 $D=0
M1300 417 75 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=15740 $D=0
M1301 418 75 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=20370 $D=0
M1302 419 415 219 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=15740 $D=0
M1303 420 416 220 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=20370 $D=0
M1304 9 419 733 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=15740 $D=0
M1305 9 420 734 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=20370 $D=0
M1306 421 733 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=15740 $D=0
M1307 422 734 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=20370 $D=0
M1308 419 74 421 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=15740 $D=0
M1309 420 74 422 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=20370 $D=0
M1310 421 417 229 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=15740 $D=0
M1311 422 418 230 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=20370 $D=0
M1312 233 423 421 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=15740 $D=0
M1313 234 424 422 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=20370 $D=0
M1314 423 76 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=15740 $D=0
M1315 424 76 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=20370 $D=0
M1316 9 77 425 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=15740 $D=0
M1317 9 77 426 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=20370 $D=0
M1318 427 78 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=15740 $D=0
M1319 428 78 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=20370 $D=0
M1320 429 425 219 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=15740 $D=0
M1321 430 426 220 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=20370 $D=0
M1322 9 429 735 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=15740 $D=0
M1323 9 430 736 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=20370 $D=0
M1324 431 735 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=15740 $D=0
M1325 432 736 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=20370 $D=0
M1326 429 77 431 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=15740 $D=0
M1327 430 77 432 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=20370 $D=0
M1328 431 427 229 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=15740 $D=0
M1329 432 428 230 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=20370 $D=0
M1330 233 433 431 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=15740 $D=0
M1331 234 434 432 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=20370 $D=0
M1332 433 79 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=15740 $D=0
M1333 434 79 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=20370 $D=0
M1334 9 80 435 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=15740 $D=0
M1335 9 80 436 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=20370 $D=0
M1336 437 81 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=15740 $D=0
M1337 438 81 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=20370 $D=0
M1338 439 435 219 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=15740 $D=0
M1339 440 436 220 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=20370 $D=0
M1340 9 439 737 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=15740 $D=0
M1341 9 440 738 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=20370 $D=0
M1342 441 737 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=15740 $D=0
M1343 442 738 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=20370 $D=0
M1344 439 80 441 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=15740 $D=0
M1345 440 80 442 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=20370 $D=0
M1346 441 437 229 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=15740 $D=0
M1347 442 438 230 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=20370 $D=0
M1348 233 443 441 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=15740 $D=0
M1349 234 444 442 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=20370 $D=0
M1350 443 82 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=15740 $D=0
M1351 444 82 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=20370 $D=0
M1352 9 83 445 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=15740 $D=0
M1353 9 83 446 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=20370 $D=0
M1354 447 84 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=15740 $D=0
M1355 448 84 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=20370 $D=0
M1356 449 445 219 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=15740 $D=0
M1357 450 446 220 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=20370 $D=0
M1358 9 449 739 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=15740 $D=0
M1359 9 450 740 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=20370 $D=0
M1360 451 739 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=15740 $D=0
M1361 452 740 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=20370 $D=0
M1362 449 83 451 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=15740 $D=0
M1363 450 83 452 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=20370 $D=0
M1364 451 447 229 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=15740 $D=0
M1365 452 448 230 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=20370 $D=0
M1366 233 453 451 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=15740 $D=0
M1367 234 454 452 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=20370 $D=0
M1368 453 85 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=15740 $D=0
M1369 454 85 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=20370 $D=0
M1370 9 86 455 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=15740 $D=0
M1371 9 86 456 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=20370 $D=0
M1372 457 87 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=15740 $D=0
M1373 458 87 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=20370 $D=0
M1374 459 455 219 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=15740 $D=0
M1375 460 456 220 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=20370 $D=0
M1376 9 459 741 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=15740 $D=0
M1377 9 460 742 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=20370 $D=0
M1378 461 741 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=15740 $D=0
M1379 462 742 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=20370 $D=0
M1380 459 86 461 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=15740 $D=0
M1381 460 86 462 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=20370 $D=0
M1382 461 457 229 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=15740 $D=0
M1383 462 458 230 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=20370 $D=0
M1384 233 463 461 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=15740 $D=0
M1385 234 464 462 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=20370 $D=0
M1386 463 88 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=15740 $D=0
M1387 464 88 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=20370 $D=0
M1388 9 89 465 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=15740 $D=0
M1389 9 89 466 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=20370 $D=0
M1390 467 90 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=15740 $D=0
M1391 468 90 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=20370 $D=0
M1392 469 465 219 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=15740 $D=0
M1393 470 466 220 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=20370 $D=0
M1394 9 469 743 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=15740 $D=0
M1395 9 470 744 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=20370 $D=0
M1396 471 743 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=15740 $D=0
M1397 472 744 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=20370 $D=0
M1398 469 89 471 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=15740 $D=0
M1399 470 89 472 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=20370 $D=0
M1400 471 467 229 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=15740 $D=0
M1401 472 468 230 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=20370 $D=0
M1402 233 473 471 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=15740 $D=0
M1403 234 474 472 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=20370 $D=0
M1404 473 91 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=15740 $D=0
M1405 474 91 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=20370 $D=0
M1406 9 92 475 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=15740 $D=0
M1407 9 92 476 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=20370 $D=0
M1408 477 93 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=15740 $D=0
M1409 478 93 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=20370 $D=0
M1410 479 475 219 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=15740 $D=0
M1411 480 476 220 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=20370 $D=0
M1412 9 479 745 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=15740 $D=0
M1413 9 480 746 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=20370 $D=0
M1414 481 745 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=15740 $D=0
M1415 482 746 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=20370 $D=0
M1416 479 92 481 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=15740 $D=0
M1417 480 92 482 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=20370 $D=0
M1418 481 477 229 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=15740 $D=0
M1419 482 478 230 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=20370 $D=0
M1420 233 483 481 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=15740 $D=0
M1421 234 484 482 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=20370 $D=0
M1422 483 94 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=15740 $D=0
M1423 484 94 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=20370 $D=0
M1424 9 95 485 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=15740 $D=0
M1425 9 95 486 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=20370 $D=0
M1426 487 96 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=15740 $D=0
M1427 488 96 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=20370 $D=0
M1428 489 485 219 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=15740 $D=0
M1429 490 486 220 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=20370 $D=0
M1430 9 489 747 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=15740 $D=0
M1431 9 490 748 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=20370 $D=0
M1432 491 747 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=15740 $D=0
M1433 492 748 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=20370 $D=0
M1434 489 95 491 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=15740 $D=0
M1435 490 95 492 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=20370 $D=0
M1436 491 487 229 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=15740 $D=0
M1437 492 488 230 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=20370 $D=0
M1438 233 493 491 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=15740 $D=0
M1439 234 494 492 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=20370 $D=0
M1440 493 97 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=15740 $D=0
M1441 494 97 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=20370 $D=0
M1442 9 98 495 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=15740 $D=0
M1443 9 98 496 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=20370 $D=0
M1444 497 99 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=15740 $D=0
M1445 498 99 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=20370 $D=0
M1446 499 495 219 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=15740 $D=0
M1447 500 496 220 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=20370 $D=0
M1448 9 499 749 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=15740 $D=0
M1449 9 500 750 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=20370 $D=0
M1450 501 749 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=15740 $D=0
M1451 502 750 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=20370 $D=0
M1452 499 98 501 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=15740 $D=0
M1453 500 98 502 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=20370 $D=0
M1454 501 497 229 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=15740 $D=0
M1455 502 498 230 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=20370 $D=0
M1456 233 503 501 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=15740 $D=0
M1457 234 504 502 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=20370 $D=0
M1458 503 100 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=15740 $D=0
M1459 504 100 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=20370 $D=0
M1460 9 101 505 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=15740 $D=0
M1461 9 101 506 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=20370 $D=0
M1462 507 102 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=15740 $D=0
M1463 508 102 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=20370 $D=0
M1464 509 505 219 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=15740 $D=0
M1465 510 506 220 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=20370 $D=0
M1466 9 509 751 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=15740 $D=0
M1467 9 510 752 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=20370 $D=0
M1468 511 751 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=15740 $D=0
M1469 512 752 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=20370 $D=0
M1470 509 101 511 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=15740 $D=0
M1471 510 101 512 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=20370 $D=0
M1472 511 507 229 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=15740 $D=0
M1473 512 508 230 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=20370 $D=0
M1474 233 513 511 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=15740 $D=0
M1475 234 514 512 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=20370 $D=0
M1476 513 103 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=15740 $D=0
M1477 514 103 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=20370 $D=0
M1478 9 104 515 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=15740 $D=0
M1479 9 104 516 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=20370 $D=0
M1480 517 105 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=15740 $D=0
M1481 518 105 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=20370 $D=0
M1482 519 515 219 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=15740 $D=0
M1483 520 516 220 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=20370 $D=0
M1484 9 519 753 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=15740 $D=0
M1485 9 520 754 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=20370 $D=0
M1486 521 753 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=15740 $D=0
M1487 522 754 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=20370 $D=0
M1488 519 104 521 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=15740 $D=0
M1489 520 104 522 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=20370 $D=0
M1490 521 517 229 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=15740 $D=0
M1491 522 518 230 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=20370 $D=0
M1492 233 523 521 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=15740 $D=0
M1493 234 524 522 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=20370 $D=0
M1494 523 107 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=15740 $D=0
M1495 524 107 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=20370 $D=0
M1496 9 109 525 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=15740 $D=0
M1497 9 109 526 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=20370 $D=0
M1498 527 110 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=15740 $D=0
M1499 528 110 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=20370 $D=0
M1500 529 525 219 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=15740 $D=0
M1501 530 526 220 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=20370 $D=0
M1502 9 529 755 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=15740 $D=0
M1503 9 530 756 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=20370 $D=0
M1504 531 755 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=15740 $D=0
M1505 532 756 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=20370 $D=0
M1506 529 109 531 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=15740 $D=0
M1507 530 109 532 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=20370 $D=0
M1508 531 527 229 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=15740 $D=0
M1509 532 528 230 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=20370 $D=0
M1510 233 533 531 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=15740 $D=0
M1511 234 534 532 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=20370 $D=0
M1512 533 113 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=15740 $D=0
M1513 534 113 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=20370 $D=0
M1514 9 114 535 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=15740 $D=0
M1515 9 114 536 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=20370 $D=0
M1516 537 115 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=15740 $D=0
M1517 538 115 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=20370 $D=0
M1518 6 537 229 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=15740 $D=0
M1519 6 538 230 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=20370 $D=0
M1520 233 535 6 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=15740 $D=0
M1521 234 536 6 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=20370 $D=0
M1522 9 541 539 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=15740 $D=0
M1523 9 542 540 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=20370 $D=0
M1524 541 116 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=15740 $D=0
M1525 542 116 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=20370 $D=0
M1526 757 229 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=15740 $D=0
M1527 758 230 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=20370 $D=0
M1528 543 541 757 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=15740 $D=0
M1529 544 542 758 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=20370 $D=0
M1530 9 543 545 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=15740 $D=0
M1531 9 544 546 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=20370 $D=0
M1532 759 545 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=15740 $D=0
M1533 760 546 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=20370 $D=0
M1534 543 539 759 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=15740 $D=0
M1535 544 540 760 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=20370 $D=0
M1536 9 549 547 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=15740 $D=0
M1537 9 550 548 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=20370 $D=0
M1538 549 116 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=15740 $D=0
M1539 550 116 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=20370 $D=0
M1540 761 233 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=15740 $D=0
M1541 762 234 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=20370 $D=0
M1542 551 549 761 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=15740 $D=0
M1543 552 550 762 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=20370 $D=0
M1544 9 551 117 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=15740 $D=0
M1545 9 552 118 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=20370 $D=0
M1546 763 117 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=15740 $D=0
M1547 764 118 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=20370 $D=0
M1548 551 547 763 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=15740 $D=0
M1549 552 548 764 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=20370 $D=0
M1550 553 119 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=15740 $D=0
M1551 554 119 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=20370 $D=0
M1552 555 119 545 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=15740 $D=0
M1553 556 119 546 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=20370 $D=0
M1554 120 553 555 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=15740 $D=0
M1555 121 554 556 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=20370 $D=0
M1556 557 122 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=15740 $D=0
M1557 558 122 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=20370 $D=0
M1558 559 122 117 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=15740 $D=0
M1559 560 122 118 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=20370 $D=0
M1560 765 557 559 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=15740 $D=0
M1561 766 558 560 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=20370 $D=0
M1562 9 117 765 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=15740 $D=0
M1563 9 118 766 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=20370 $D=0
M1564 561 123 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=15740 $D=0
M1565 562 123 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=20370 $D=0
M1566 563 123 559 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=15740 $D=0
M1567 564 123 560 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=20370 $D=0
M1568 11 561 563 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=15740 $D=0
M1569 12 562 564 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=20370 $D=0
M1570 566 565 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=15740 $D=0
M1571 567 124 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=20370 $D=0
M1572 9 570 568 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=15740 $D=0
M1573 9 571 569 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=20370 $D=0
M1574 572 555 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=15740 $D=0
M1575 573 556 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=20370 $D=0
M1576 570 555 565 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=15740 $D=0
M1577 571 556 124 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=20370 $D=0
M1578 566 572 570 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=15740 $D=0
M1579 567 573 571 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=20370 $D=0
M1580 574 568 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=15740 $D=0
M1581 575 569 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=20370 $D=0
M1582 125 568 563 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=15740 $D=0
M1583 565 569 564 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=20370 $D=0
M1584 555 574 125 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=15740 $D=0
M1585 556 575 565 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=20370 $D=0
M1586 576 125 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=15740 $D=0
M1587 577 565 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=20370 $D=0
M1588 578 568 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=15740 $D=0
M1589 579 569 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=20370 $D=0
M1590 580 568 576 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=15740 $D=0
M1591 581 569 577 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=20370 $D=0
M1592 563 578 580 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=15740 $D=0
M1593 564 579 581 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=20370 $D=0
M1594 777 555 9 9 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=15380 $D=0
M1595 778 556 9 9 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=20010 $D=0
M1596 582 563 777 9 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=15380 $D=0
M1597 583 564 778 9 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=20010 $D=0
M1598 584 580 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=15740 $D=0
M1599 585 581 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=20370 $D=0
M1600 586 555 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=15740 $D=0
M1601 587 556 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=20370 $D=0
M1602 9 563 586 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=15740 $D=0
M1603 9 564 587 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=20370 $D=0
M1604 588 555 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=15740 $D=0
M1605 589 556 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=20370 $D=0
M1606 9 563 588 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=15740 $D=0
M1607 9 564 589 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=20370 $D=0
M1608 779 555 9 9 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=15560 $D=0
M1609 780 556 9 9 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=20190 $D=0
M1610 592 563 779 9 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=15560 $D=0
M1611 593 564 780 9 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=20190 $D=0
M1612 9 588 592 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=15740 $D=0
M1613 9 589 593 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=20370 $D=0
M1614 594 128 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=15740 $D=0
M1615 595 128 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=20370 $D=0
M1616 596 128 582 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=15740 $D=0
M1617 597 128 583 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=20370 $D=0
M1618 586 594 596 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=15740 $D=0
M1619 587 595 597 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=20370 $D=0
M1620 598 128 584 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=15740 $D=0
M1621 599 128 585 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=20370 $D=0
M1622 592 594 598 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=15740 $D=0
M1623 593 595 599 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=20370 $D=0
M1624 600 129 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=15740 $D=0
M1625 601 129 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=20370 $D=0
M1626 602 129 598 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=15740 $D=0
M1627 603 129 599 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=20370 $D=0
M1628 596 600 602 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=15740 $D=0
M1629 597 601 603 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=20370 $D=0
M1630 13 602 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=15740 $D=0
M1631 14 603 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=20370 $D=0
M1632 604 130 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=15740 $D=0
M1633 605 130 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=20370 $D=0
M1634 606 130 131 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=15740 $D=0
M1635 607 130 132 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=20370 $D=0
M1636 133 604 606 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=15740 $D=0
M1637 134 605 607 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=20370 $D=0
M1638 608 130 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=15740 $D=0
M1639 609 130 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=20370 $D=0
M1640 610 130 135 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=15740 $D=0
M1641 611 130 136 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=20370 $D=0
M1642 137 608 610 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=15740 $D=0
M1643 138 609 611 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=20370 $D=0
M1644 612 130 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=15740 $D=0
M1645 613 130 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=20370 $D=0
M1646 614 130 126 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=15740 $D=0
M1647 615 130 127 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=20370 $D=0
M1648 139 612 614 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=15740 $D=0
M1649 140 613 615 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=20370 $D=0
M1650 616 130 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=15740 $D=0
M1651 617 130 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=20370 $D=0
M1652 618 130 142 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=15740 $D=0
M1653 619 130 143 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=20370 $D=0
M1654 139 616 618 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=15740 $D=0
M1655 139 617 619 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=20370 $D=0
M1656 620 130 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=15740 $D=0
M1657 621 130 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=20370 $D=0
M1658 622 130 144 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=15740 $D=0
M1659 623 130 145 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=20370 $D=0
M1660 139 620 622 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=15740 $D=0
M1661 139 621 623 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=20370 $D=0
M1662 9 555 767 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=15740 $D=0
M1663 9 556 768 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=20370 $D=0
M1664 134 767 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=15740 $D=0
M1665 131 768 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=20370 $D=0
M1666 624 146 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=15740 $D=0
M1667 625 146 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=20370 $D=0
M1668 147 146 134 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=15740 $D=0
M1669 148 146 131 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=20370 $D=0
M1670 606 624 147 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=15740 $D=0
M1671 607 625 148 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=20370 $D=0
M1672 626 149 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=15740 $D=0
M1673 627 149 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=20370 $D=0
M1674 150 149 147 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=15740 $D=0
M1675 106 149 148 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=20370 $D=0
M1676 610 626 150 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=15740 $D=0
M1677 611 627 106 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=20370 $D=0
M1678 628 151 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=15740 $D=0
M1679 629 151 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=20370 $D=0
M1680 152 151 150 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=15740 $D=0
M1681 111 151 106 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=20370 $D=0
M1682 614 628 152 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=15740 $D=0
M1683 615 629 111 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=20370 $D=0
M1684 630 153 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=15740 $D=0
M1685 631 153 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=20370 $D=0
M1686 154 153 152 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=15740 $D=0
M1687 155 153 111 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=20370 $D=0
M1688 618 630 154 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=15740 $D=0
M1689 619 631 155 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=20370 $D=0
M1690 632 156 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=15740 $D=0
M1691 633 156 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=20370 $D=0
M1692 205 156 154 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=15740 $D=0
M1693 206 156 155 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=20370 $D=0
M1694 622 632 205 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=15740 $D=0
M1695 623 633 206 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=20370 $D=0
M1696 634 157 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=15740 $D=0
M1697 635 157 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=20370 $D=0
M1698 636 157 117 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=15740 $D=0
M1699 637 157 118 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=20370 $D=0
M1700 11 634 636 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=15740 $D=0
M1701 12 635 637 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=20370 $D=0
M1702 638 545 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=15740 $D=0
M1703 639 546 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=20370 $D=0
M1704 9 636 638 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=15740 $D=0
M1705 9 637 639 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=20370 $D=0
M1706 781 545 9 9 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=15560 $D=0
M1707 782 546 9 9 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=20190 $D=0
M1708 642 636 781 9 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=15560 $D=0
M1709 643 637 782 9 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=20190 $D=0
M1710 9 638 642 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=15740 $D=0
M1711 9 639 643 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=20370 $D=0
M1712 769 158 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=15740 $D=0
M1713 770 644 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=20370 $D=0
M1714 9 642 769 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=15740 $D=0
M1715 9 643 770 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=20370 $D=0
M1716 644 769 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=15740 $D=0
M1717 159 770 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=20370 $D=0
M1718 783 545 9 9 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=15380 $D=0
M1719 784 546 9 9 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=20010 $D=0
M1720 645 647 783 9 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=15380 $D=0
M1721 646 648 784 9 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=20010 $D=0
M1722 647 636 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=15740 $D=0
M1723 648 637 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=20370 $D=0
M1724 649 645 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=15740 $D=0
M1725 650 646 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=20370 $D=0
M1726 9 158 649 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=15740 $D=0
M1727 9 644 650 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=20370 $D=0
M1728 652 160 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=15740 $D=0
M1729 653 651 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=20370 $D=0
M1730 651 649 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=15740 $D=0
M1731 161 650 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=20370 $D=0
M1732 9 652 651 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=15740 $D=0
M1733 9 653 161 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=20370 $D=0
M1734 655 654 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=15740 $D=0
M1735 656 162 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=20370 $D=0
M1736 9 659 657 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=15740 $D=0
M1737 9 660 658 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=20370 $D=0
M1738 661 120 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=15740 $D=0
M1739 662 121 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=20370 $D=0
M1740 659 120 654 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=15740 $D=0
M1741 660 121 162 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=20370 $D=0
M1742 655 661 659 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=15740 $D=0
M1743 656 662 660 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=20370 $D=0
M1744 663 657 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=15740 $D=0
M1745 664 658 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=20370 $D=0
M1746 163 657 6 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=15740 $D=0
M1747 654 658 6 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=20370 $D=0
M1748 120 663 163 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=15740 $D=0
M1749 121 664 654 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=20370 $D=0
M1750 665 163 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=15740 $D=0
M1751 666 654 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=20370 $D=0
M1752 667 657 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=15740 $D=0
M1753 668 658 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=20370 $D=0
M1754 207 657 665 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=15740 $D=0
M1755 208 658 666 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=20370 $D=0
M1756 6 667 207 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=15740 $D=0
M1757 6 668 208 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=20370 $D=0
M1758 669 164 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=15740 $D=0
M1759 670 164 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=20370 $D=0
M1760 671 164 207 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=15740 $D=0
M1761 672 164 208 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=20370 $D=0
M1762 13 669 671 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=15740 $D=0
M1763 14 670 672 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=20370 $D=0
M1764 673 165 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=15740 $D=0
M1765 674 165 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=20370 $D=0
M1766 675 165 671 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=15740 $D=0
M1767 676 165 672 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=20370 $D=0
M1768 6 673 675 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=15740 $D=0
M1769 6 674 676 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=20370 $D=0
M1770 677 116 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=15740 $D=0
M1771 678 116 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=20370 $D=0
M1772 9 677 679 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=15740 $D=0
M1773 9 678 680 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=20370 $D=0
M1774 681 116 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=15740 $D=0
M1775 682 116 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=20370 $D=0
M1776 683 679 675 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=15740 $D=0
M1777 684 680 676 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=20370 $D=0
M1778 9 683 771 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=15740 $D=0
M1779 9 684 772 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=20370 $D=0
M1780 685 771 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=15740 $D=0
M1781 686 772 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=20370 $D=0
M1782 683 677 685 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=15740 $D=0
M1783 684 678 686 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=20370 $D=0
M1784 687 681 685 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=15740 $D=0
M1785 688 682 686 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=20370 $D=0
M1786 9 691 689 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=15740 $D=0
M1787 9 692 690 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=20370 $D=0
M1788 691 116 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=15740 $D=0
M1789 692 116 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=20370 $D=0
M1790 773 687 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=15740 $D=0
M1791 774 688 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=20370 $D=0
M1792 693 691 773 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=15740 $D=0
M1793 694 692 774 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=20370 $D=0
M1794 9 693 120 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=15740 $D=0
M1795 9 694 121 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=20370 $D=0
M1796 775 120 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=15740 $D=0
M1797 776 121 9 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=20370 $D=0
M1798 693 689 775 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=15740 $D=0
M1799 694 690 776 9 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=20370 $D=0
.ENDS
***************************************
.SUBCKT ICV_41 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 116 117 118 119 120 121
+ 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141
+ 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161
+ 162 163 164 165 166 167
** N=1097 EP=166 IP=2241 FDC=2700
M0 169 1 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=600 $D=1
M1 170 1 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=5230 $D=1
M2 171 1 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=9860 $D=1
M3 172 169 2 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=600 $D=1
M4 173 170 3 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=5230 $D=1
M5 174 171 4 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=9860 $D=1
M6 7 1 172 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=600 $D=1
M7 7 1 173 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=5230 $D=1
M8 7 1 174 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=9860 $D=1
M9 175 169 5 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=600 $D=1
M10 176 170 5 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=5230 $D=1
M11 177 171 5 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=9860 $D=1
M12 6 1 175 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=600 $D=1
M13 6 1 176 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=5230 $D=1
M14 6 1 177 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=9860 $D=1
M15 178 169 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=600 $D=1
M16 179 170 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=5230 $D=1
M17 180 171 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=9860 $D=1
M18 7 1 178 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=600 $D=1
M19 7 1 179 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=5230 $D=1
M20 7 1 180 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=9860 $D=1
M21 184 181 178 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=600 $D=1
M22 185 182 179 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=5230 $D=1
M23 186 183 180 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=9860 $D=1
M24 181 8 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=600 $D=1
M25 182 8 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=5230 $D=1
M26 183 8 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=9860 $D=1
M27 187 181 175 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=600 $D=1
M28 188 182 176 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=5230 $D=1
M29 189 183 177 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=9860 $D=1
M30 172 8 187 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=600 $D=1
M31 173 8 188 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=5230 $D=1
M32 174 8 189 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=9860 $D=1
M33 190 9 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=600 $D=1
M34 191 9 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=5230 $D=1
M35 192 9 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=9860 $D=1
M36 193 190 187 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=600 $D=1
M37 194 191 188 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=5230 $D=1
M38 195 192 189 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=9860 $D=1
M39 184 9 193 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=600 $D=1
M40 185 9 194 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=5230 $D=1
M41 186 9 195 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=9860 $D=1
M42 196 11 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=600 $D=1
M43 197 11 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=5230 $D=1
M44 198 11 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=9860 $D=1
M45 199 196 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=600 $D=1
M46 200 197 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=5230 $D=1
M47 201 198 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=9860 $D=1
M48 12 11 199 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=600 $D=1
M49 13 11 200 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=5230 $D=1
M50 14 11 201 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=9860 $D=1
M51 202 196 15 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=600 $D=1
M52 203 197 16 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=5230 $D=1
M53 204 198 17 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=9860 $D=1
M54 205 11 202 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=600 $D=1
M55 206 11 203 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=5230 $D=1
M56 207 11 204 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=9860 $D=1
M57 211 196 208 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=600 $D=1
M58 212 197 209 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=5230 $D=1
M59 213 198 210 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=9860 $D=1
M60 193 11 211 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=600 $D=1
M61 194 11 212 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=5230 $D=1
M62 195 11 213 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=9860 $D=1
M63 217 214 211 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=600 $D=1
M64 218 215 212 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=5230 $D=1
M65 219 216 213 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=9860 $D=1
M66 214 18 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=600 $D=1
M67 215 18 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=5230 $D=1
M68 216 18 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=9860 $D=1
M69 220 214 202 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=600 $D=1
M70 221 215 203 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=5230 $D=1
M71 222 216 204 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=9860 $D=1
M72 199 18 220 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=600 $D=1
M73 200 18 221 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=5230 $D=1
M74 201 18 222 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=9860 $D=1
M75 223 19 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=600 $D=1
M76 224 19 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=5230 $D=1
M77 225 19 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=9860 $D=1
M78 226 223 220 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=600 $D=1
M79 227 224 221 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=5230 $D=1
M80 228 225 222 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=9860 $D=1
M81 217 19 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=600 $D=1
M82 218 19 227 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=5230 $D=1
M83 219 19 228 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=9860 $D=1
M84 7 20 229 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=600 $D=1
M85 7 20 230 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=5230 $D=1
M86 7 20 231 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=9860 $D=1
M87 232 21 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=600 $D=1
M88 233 21 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=5230 $D=1
M89 234 21 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=9860 $D=1
M90 235 20 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=600 $D=1
M91 236 20 227 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=5230 $D=1
M92 237 20 228 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=9860 $D=1
M93 7 235 945 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=600 $D=1
M94 7 236 946 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=5230 $D=1
M95 7 237 947 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=9860 $D=1
M96 238 945 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=600 $D=1
M97 239 946 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=5230 $D=1
M98 240 947 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=9860 $D=1
M99 235 229 238 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=600 $D=1
M100 236 230 239 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=5230 $D=1
M101 237 231 240 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=9860 $D=1
M102 238 21 241 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=600 $D=1
M103 239 21 242 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=5230 $D=1
M104 240 21 243 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=9860 $D=1
M105 247 22 238 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=600 $D=1
M106 248 22 239 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=5230 $D=1
M107 249 22 240 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=9860 $D=1
M108 244 22 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=600 $D=1
M109 245 22 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=5230 $D=1
M110 246 22 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=9860 $D=1
M111 7 23 250 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=600 $D=1
M112 7 23 251 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=5230 $D=1
M113 7 23 252 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=9860 $D=1
M114 253 24 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=600 $D=1
M115 254 24 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=5230 $D=1
M116 255 24 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=9860 $D=1
M117 256 23 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=600 $D=1
M118 257 23 227 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=5230 $D=1
M119 258 23 228 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=9860 $D=1
M120 7 256 948 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=600 $D=1
M121 7 257 949 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=5230 $D=1
M122 7 258 950 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=9860 $D=1
M123 259 948 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=600 $D=1
M124 260 949 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=5230 $D=1
M125 261 950 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=9860 $D=1
M126 256 250 259 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=600 $D=1
M127 257 251 260 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=5230 $D=1
M128 258 252 261 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=9860 $D=1
M129 259 24 241 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=600 $D=1
M130 260 24 242 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=5230 $D=1
M131 261 24 243 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=9860 $D=1
M132 247 25 259 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=600 $D=1
M133 248 25 260 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=5230 $D=1
M134 249 25 261 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=9860 $D=1
M135 262 25 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=600 $D=1
M136 263 25 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=5230 $D=1
M137 264 25 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=9860 $D=1
M138 7 26 265 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=600 $D=1
M139 7 26 266 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=5230 $D=1
M140 7 26 267 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=9860 $D=1
M141 268 27 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=600 $D=1
M142 269 27 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=5230 $D=1
M143 270 27 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=9860 $D=1
M144 271 26 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=600 $D=1
M145 272 26 227 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=5230 $D=1
M146 273 26 228 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=9860 $D=1
M147 7 271 951 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=600 $D=1
M148 7 272 952 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=5230 $D=1
M149 7 273 953 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=9860 $D=1
M150 274 951 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=600 $D=1
M151 275 952 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=5230 $D=1
M152 276 953 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=9860 $D=1
M153 271 265 274 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=600 $D=1
M154 272 266 275 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=5230 $D=1
M155 273 267 276 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=9860 $D=1
M156 274 27 241 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=600 $D=1
M157 275 27 242 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=5230 $D=1
M158 276 27 243 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=9860 $D=1
M159 247 28 274 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=600 $D=1
M160 248 28 275 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=5230 $D=1
M161 249 28 276 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=9860 $D=1
M162 277 28 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=600 $D=1
M163 278 28 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=5230 $D=1
M164 279 28 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=9860 $D=1
M165 7 29 280 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=600 $D=1
M166 7 29 281 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=5230 $D=1
M167 7 29 282 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=9860 $D=1
M168 283 30 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=600 $D=1
M169 284 30 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=5230 $D=1
M170 285 30 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=9860 $D=1
M171 286 29 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=600 $D=1
M172 287 29 227 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=5230 $D=1
M173 288 29 228 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=9860 $D=1
M174 7 286 954 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=600 $D=1
M175 7 287 955 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=5230 $D=1
M176 7 288 956 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=9860 $D=1
M177 289 954 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=600 $D=1
M178 290 955 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=5230 $D=1
M179 291 956 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=9860 $D=1
M180 286 280 289 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=600 $D=1
M181 287 281 290 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=5230 $D=1
M182 288 282 291 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=9860 $D=1
M183 289 30 241 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=600 $D=1
M184 290 30 242 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=5230 $D=1
M185 291 30 243 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=9860 $D=1
M186 247 31 289 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=600 $D=1
M187 248 31 290 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=5230 $D=1
M188 249 31 291 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=9860 $D=1
M189 292 31 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=600 $D=1
M190 293 31 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=5230 $D=1
M191 294 31 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=9860 $D=1
M192 7 32 295 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=600 $D=1
M193 7 32 296 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=5230 $D=1
M194 7 32 297 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=9860 $D=1
M195 298 33 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=600 $D=1
M196 299 33 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=5230 $D=1
M197 300 33 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=9860 $D=1
M198 301 32 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=600 $D=1
M199 302 32 227 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=5230 $D=1
M200 303 32 228 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=9860 $D=1
M201 7 301 957 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=600 $D=1
M202 7 302 958 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=5230 $D=1
M203 7 303 959 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=9860 $D=1
M204 304 957 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=600 $D=1
M205 305 958 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=5230 $D=1
M206 306 959 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=9860 $D=1
M207 301 295 304 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=600 $D=1
M208 302 296 305 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=5230 $D=1
M209 303 297 306 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=9860 $D=1
M210 304 33 241 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=600 $D=1
M211 305 33 242 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=5230 $D=1
M212 306 33 243 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=9860 $D=1
M213 247 34 304 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=600 $D=1
M214 248 34 305 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=5230 $D=1
M215 249 34 306 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=9860 $D=1
M216 307 34 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=600 $D=1
M217 308 34 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=5230 $D=1
M218 309 34 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=9860 $D=1
M219 7 35 310 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=600 $D=1
M220 7 35 311 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=5230 $D=1
M221 7 35 312 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=9860 $D=1
M222 313 36 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=600 $D=1
M223 314 36 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=5230 $D=1
M224 315 36 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=9860 $D=1
M225 316 35 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=600 $D=1
M226 317 35 227 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=5230 $D=1
M227 318 35 228 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=9860 $D=1
M228 7 316 960 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=600 $D=1
M229 7 317 961 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=5230 $D=1
M230 7 318 962 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=9860 $D=1
M231 319 960 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=600 $D=1
M232 320 961 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=5230 $D=1
M233 321 962 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=9860 $D=1
M234 316 310 319 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=600 $D=1
M235 317 311 320 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=5230 $D=1
M236 318 312 321 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=9860 $D=1
M237 319 36 241 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=600 $D=1
M238 320 36 242 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=5230 $D=1
M239 321 36 243 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=9860 $D=1
M240 247 37 319 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=600 $D=1
M241 248 37 320 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=5230 $D=1
M242 249 37 321 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=9860 $D=1
M243 322 37 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=600 $D=1
M244 323 37 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=5230 $D=1
M245 324 37 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=9860 $D=1
M246 7 38 325 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=600 $D=1
M247 7 38 326 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=5230 $D=1
M248 7 38 327 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=9860 $D=1
M249 328 39 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=600 $D=1
M250 329 39 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=5230 $D=1
M251 330 39 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=9860 $D=1
M252 331 38 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=600 $D=1
M253 332 38 227 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=5230 $D=1
M254 333 38 228 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=9860 $D=1
M255 7 331 963 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=600 $D=1
M256 7 332 964 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=5230 $D=1
M257 7 333 965 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=9860 $D=1
M258 334 963 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=600 $D=1
M259 335 964 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=5230 $D=1
M260 336 965 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=9860 $D=1
M261 331 325 334 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=600 $D=1
M262 332 326 335 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=5230 $D=1
M263 333 327 336 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=9860 $D=1
M264 334 39 241 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=600 $D=1
M265 335 39 242 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=5230 $D=1
M266 336 39 243 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=9860 $D=1
M267 247 40 334 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=600 $D=1
M268 248 40 335 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=5230 $D=1
M269 249 40 336 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=9860 $D=1
M270 337 40 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=600 $D=1
M271 338 40 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=5230 $D=1
M272 339 40 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=9860 $D=1
M273 7 41 340 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=600 $D=1
M274 7 41 341 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=5230 $D=1
M275 7 41 342 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=9860 $D=1
M276 343 42 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=600 $D=1
M277 344 42 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=5230 $D=1
M278 345 42 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=9860 $D=1
M279 346 41 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=600 $D=1
M280 347 41 227 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=5230 $D=1
M281 348 41 228 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=9860 $D=1
M282 7 346 966 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=600 $D=1
M283 7 347 967 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=5230 $D=1
M284 7 348 968 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=9860 $D=1
M285 349 966 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=600 $D=1
M286 350 967 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=5230 $D=1
M287 351 968 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=9860 $D=1
M288 346 340 349 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=600 $D=1
M289 347 341 350 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=5230 $D=1
M290 348 342 351 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=9860 $D=1
M291 349 42 241 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=600 $D=1
M292 350 42 242 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=5230 $D=1
M293 351 42 243 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=9860 $D=1
M294 247 43 349 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=600 $D=1
M295 248 43 350 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=5230 $D=1
M296 249 43 351 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=9860 $D=1
M297 352 43 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=600 $D=1
M298 353 43 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=5230 $D=1
M299 354 43 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=9860 $D=1
M300 7 44 355 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=600 $D=1
M301 7 44 356 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=5230 $D=1
M302 7 44 357 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=9860 $D=1
M303 358 45 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=600 $D=1
M304 359 45 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=5230 $D=1
M305 360 45 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=9860 $D=1
M306 361 44 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=600 $D=1
M307 362 44 227 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=5230 $D=1
M308 363 44 228 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=9860 $D=1
M309 7 361 969 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=600 $D=1
M310 7 362 970 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=5230 $D=1
M311 7 363 971 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=9860 $D=1
M312 364 969 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=600 $D=1
M313 365 970 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=5230 $D=1
M314 366 971 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=9860 $D=1
M315 361 355 364 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=600 $D=1
M316 362 356 365 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=5230 $D=1
M317 363 357 366 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=9860 $D=1
M318 364 45 241 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=600 $D=1
M319 365 45 242 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=5230 $D=1
M320 366 45 243 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=9860 $D=1
M321 247 46 364 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=600 $D=1
M322 248 46 365 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=5230 $D=1
M323 249 46 366 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=9860 $D=1
M324 367 46 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=600 $D=1
M325 368 46 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=5230 $D=1
M326 369 46 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=9860 $D=1
M327 7 47 370 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=600 $D=1
M328 7 47 371 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=5230 $D=1
M329 7 47 372 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=9860 $D=1
M330 373 48 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=600 $D=1
M331 374 48 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=5230 $D=1
M332 375 48 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=9860 $D=1
M333 376 47 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=600 $D=1
M334 377 47 227 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=5230 $D=1
M335 378 47 228 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=9860 $D=1
M336 7 376 972 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=600 $D=1
M337 7 377 973 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=5230 $D=1
M338 7 378 974 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=9860 $D=1
M339 379 972 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=600 $D=1
M340 380 973 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=5230 $D=1
M341 381 974 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=9860 $D=1
M342 376 370 379 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=600 $D=1
M343 377 371 380 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=5230 $D=1
M344 378 372 381 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=9860 $D=1
M345 379 48 241 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=600 $D=1
M346 380 48 242 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=5230 $D=1
M347 381 48 243 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=9860 $D=1
M348 247 49 379 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=600 $D=1
M349 248 49 380 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=5230 $D=1
M350 249 49 381 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=9860 $D=1
M351 382 49 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=600 $D=1
M352 383 49 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=5230 $D=1
M353 384 49 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=9860 $D=1
M354 7 50 385 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=600 $D=1
M355 7 50 386 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=5230 $D=1
M356 7 50 387 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=9860 $D=1
M357 388 51 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=600 $D=1
M358 389 51 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=5230 $D=1
M359 390 51 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=9860 $D=1
M360 391 50 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=600 $D=1
M361 392 50 227 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=5230 $D=1
M362 393 50 228 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=9860 $D=1
M363 7 391 975 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=600 $D=1
M364 7 392 976 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=5230 $D=1
M365 7 393 977 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=9860 $D=1
M366 394 975 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=600 $D=1
M367 395 976 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=5230 $D=1
M368 396 977 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=9860 $D=1
M369 391 385 394 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=600 $D=1
M370 392 386 395 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=5230 $D=1
M371 393 387 396 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=9860 $D=1
M372 394 51 241 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=600 $D=1
M373 395 51 242 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=5230 $D=1
M374 396 51 243 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=9860 $D=1
M375 247 52 394 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=600 $D=1
M376 248 52 395 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=5230 $D=1
M377 249 52 396 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=9860 $D=1
M378 397 52 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=600 $D=1
M379 398 52 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=5230 $D=1
M380 399 52 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=9860 $D=1
M381 7 53 400 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=600 $D=1
M382 7 53 401 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=5230 $D=1
M383 7 53 402 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=9860 $D=1
M384 403 54 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=600 $D=1
M385 404 54 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=5230 $D=1
M386 405 54 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=9860 $D=1
M387 406 53 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=600 $D=1
M388 407 53 227 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=5230 $D=1
M389 408 53 228 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=9860 $D=1
M390 7 406 978 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=600 $D=1
M391 7 407 979 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=5230 $D=1
M392 7 408 980 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=9860 $D=1
M393 409 978 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=600 $D=1
M394 410 979 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=5230 $D=1
M395 411 980 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=9860 $D=1
M396 406 400 409 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=600 $D=1
M397 407 401 410 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=5230 $D=1
M398 408 402 411 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=9860 $D=1
M399 409 54 241 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=600 $D=1
M400 410 54 242 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=5230 $D=1
M401 411 54 243 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=9860 $D=1
M402 247 55 409 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=600 $D=1
M403 248 55 410 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=5230 $D=1
M404 249 55 411 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=9860 $D=1
M405 412 55 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=600 $D=1
M406 413 55 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=5230 $D=1
M407 414 55 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=9860 $D=1
M408 7 56 415 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=600 $D=1
M409 7 56 416 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=5230 $D=1
M410 7 56 417 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=9860 $D=1
M411 418 57 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=600 $D=1
M412 419 57 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=5230 $D=1
M413 420 57 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=9860 $D=1
M414 421 56 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=600 $D=1
M415 422 56 227 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=5230 $D=1
M416 423 56 228 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=9860 $D=1
M417 7 421 981 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=600 $D=1
M418 7 422 982 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=5230 $D=1
M419 7 423 983 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=9860 $D=1
M420 424 981 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=600 $D=1
M421 425 982 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=5230 $D=1
M422 426 983 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=9860 $D=1
M423 421 415 424 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=600 $D=1
M424 422 416 425 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=5230 $D=1
M425 423 417 426 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=9860 $D=1
M426 424 57 241 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=600 $D=1
M427 425 57 242 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=5230 $D=1
M428 426 57 243 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=9860 $D=1
M429 247 58 424 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=600 $D=1
M430 248 58 425 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=5230 $D=1
M431 249 58 426 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=9860 $D=1
M432 427 58 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=600 $D=1
M433 428 58 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=5230 $D=1
M434 429 58 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=9860 $D=1
M435 7 59 430 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=600 $D=1
M436 7 59 431 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=5230 $D=1
M437 7 59 432 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=9860 $D=1
M438 433 60 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=600 $D=1
M439 434 60 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=5230 $D=1
M440 435 60 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=9860 $D=1
M441 436 59 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=600 $D=1
M442 437 59 227 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=5230 $D=1
M443 438 59 228 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=9860 $D=1
M444 7 436 984 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=600 $D=1
M445 7 437 985 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=5230 $D=1
M446 7 438 986 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=9860 $D=1
M447 439 984 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=600 $D=1
M448 440 985 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=5230 $D=1
M449 441 986 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=9860 $D=1
M450 436 430 439 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=600 $D=1
M451 437 431 440 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=5230 $D=1
M452 438 432 441 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=9860 $D=1
M453 439 60 241 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=600 $D=1
M454 440 60 242 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=5230 $D=1
M455 441 60 243 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=9860 $D=1
M456 247 61 439 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=600 $D=1
M457 248 61 440 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=5230 $D=1
M458 249 61 441 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=9860 $D=1
M459 442 61 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=600 $D=1
M460 443 61 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=5230 $D=1
M461 444 61 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=9860 $D=1
M462 7 62 445 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=600 $D=1
M463 7 62 446 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=5230 $D=1
M464 7 62 447 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=9860 $D=1
M465 448 63 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=600 $D=1
M466 449 63 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=5230 $D=1
M467 450 63 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=9860 $D=1
M468 451 62 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=600 $D=1
M469 452 62 227 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=5230 $D=1
M470 453 62 228 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=9860 $D=1
M471 7 451 987 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=600 $D=1
M472 7 452 988 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=5230 $D=1
M473 7 453 989 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=9860 $D=1
M474 454 987 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=600 $D=1
M475 455 988 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=5230 $D=1
M476 456 989 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=9860 $D=1
M477 451 445 454 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=600 $D=1
M478 452 446 455 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=5230 $D=1
M479 453 447 456 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=9860 $D=1
M480 454 63 241 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=600 $D=1
M481 455 63 242 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=5230 $D=1
M482 456 63 243 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=9860 $D=1
M483 247 64 454 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=600 $D=1
M484 248 64 455 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=5230 $D=1
M485 249 64 456 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=9860 $D=1
M486 457 64 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=600 $D=1
M487 458 64 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=5230 $D=1
M488 459 64 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=9860 $D=1
M489 7 65 460 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=600 $D=1
M490 7 65 461 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=5230 $D=1
M491 7 65 462 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=9860 $D=1
M492 463 66 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=600 $D=1
M493 464 66 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=5230 $D=1
M494 465 66 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=9860 $D=1
M495 466 65 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=600 $D=1
M496 467 65 227 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=5230 $D=1
M497 468 65 228 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=9860 $D=1
M498 7 466 990 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=600 $D=1
M499 7 467 991 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=5230 $D=1
M500 7 468 992 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=9860 $D=1
M501 469 990 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=600 $D=1
M502 470 991 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=5230 $D=1
M503 471 992 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=9860 $D=1
M504 466 460 469 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=600 $D=1
M505 467 461 470 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=5230 $D=1
M506 468 462 471 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=9860 $D=1
M507 469 66 241 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=600 $D=1
M508 470 66 242 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=5230 $D=1
M509 471 66 243 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=9860 $D=1
M510 247 67 469 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=600 $D=1
M511 248 67 470 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=5230 $D=1
M512 249 67 471 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=9860 $D=1
M513 472 67 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=600 $D=1
M514 473 67 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=5230 $D=1
M515 474 67 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=9860 $D=1
M516 7 68 475 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=600 $D=1
M517 7 68 476 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=5230 $D=1
M518 7 68 477 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=9860 $D=1
M519 478 69 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=600 $D=1
M520 479 69 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=5230 $D=1
M521 480 69 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=9860 $D=1
M522 481 68 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=600 $D=1
M523 482 68 227 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=5230 $D=1
M524 483 68 228 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=9860 $D=1
M525 7 481 993 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=600 $D=1
M526 7 482 994 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=5230 $D=1
M527 7 483 995 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=9860 $D=1
M528 484 993 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=600 $D=1
M529 485 994 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=5230 $D=1
M530 486 995 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=9860 $D=1
M531 481 475 484 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=600 $D=1
M532 482 476 485 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=5230 $D=1
M533 483 477 486 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=9860 $D=1
M534 484 69 241 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=600 $D=1
M535 485 69 242 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=5230 $D=1
M536 486 69 243 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=9860 $D=1
M537 247 70 484 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=600 $D=1
M538 248 70 485 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=5230 $D=1
M539 249 70 486 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=9860 $D=1
M540 487 70 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=600 $D=1
M541 488 70 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=5230 $D=1
M542 489 70 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=9860 $D=1
M543 7 71 490 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=600 $D=1
M544 7 71 491 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=5230 $D=1
M545 7 71 492 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=9860 $D=1
M546 493 72 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=600 $D=1
M547 494 72 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=5230 $D=1
M548 495 72 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=9860 $D=1
M549 496 71 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=600 $D=1
M550 497 71 227 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=5230 $D=1
M551 498 71 228 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=9860 $D=1
M552 7 496 996 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=600 $D=1
M553 7 497 997 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=5230 $D=1
M554 7 498 998 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=9860 $D=1
M555 499 996 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=600 $D=1
M556 500 997 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=5230 $D=1
M557 501 998 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=9860 $D=1
M558 496 490 499 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=600 $D=1
M559 497 491 500 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=5230 $D=1
M560 498 492 501 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=9860 $D=1
M561 499 72 241 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=600 $D=1
M562 500 72 242 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=5230 $D=1
M563 501 72 243 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=9860 $D=1
M564 247 73 499 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=600 $D=1
M565 248 73 500 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=5230 $D=1
M566 249 73 501 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=9860 $D=1
M567 502 73 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=600 $D=1
M568 503 73 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=5230 $D=1
M569 504 73 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=9860 $D=1
M570 7 74 505 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=600 $D=1
M571 7 74 506 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=5230 $D=1
M572 7 74 507 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=9860 $D=1
M573 508 75 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=600 $D=1
M574 509 75 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=5230 $D=1
M575 510 75 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=9860 $D=1
M576 511 74 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=600 $D=1
M577 512 74 227 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=5230 $D=1
M578 513 74 228 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=9860 $D=1
M579 7 511 999 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=600 $D=1
M580 7 512 1000 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=5230 $D=1
M581 7 513 1001 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=9860 $D=1
M582 514 999 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=600 $D=1
M583 515 1000 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=5230 $D=1
M584 516 1001 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=9860 $D=1
M585 511 505 514 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=600 $D=1
M586 512 506 515 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=5230 $D=1
M587 513 507 516 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=9860 $D=1
M588 514 75 241 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=600 $D=1
M589 515 75 242 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=5230 $D=1
M590 516 75 243 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=9860 $D=1
M591 247 76 514 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=600 $D=1
M592 248 76 515 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=5230 $D=1
M593 249 76 516 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=9860 $D=1
M594 517 76 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=600 $D=1
M595 518 76 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=5230 $D=1
M596 519 76 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=9860 $D=1
M597 7 77 520 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=600 $D=1
M598 7 77 521 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=5230 $D=1
M599 7 77 522 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=9860 $D=1
M600 523 78 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=600 $D=1
M601 524 78 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=5230 $D=1
M602 525 78 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=9860 $D=1
M603 526 77 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=600 $D=1
M604 527 77 227 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=5230 $D=1
M605 528 77 228 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=9860 $D=1
M606 7 526 1002 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=600 $D=1
M607 7 527 1003 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=5230 $D=1
M608 7 528 1004 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=9860 $D=1
M609 529 1002 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=600 $D=1
M610 530 1003 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=5230 $D=1
M611 531 1004 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=9860 $D=1
M612 526 520 529 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=600 $D=1
M613 527 521 530 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=5230 $D=1
M614 528 522 531 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=9860 $D=1
M615 529 78 241 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=600 $D=1
M616 530 78 242 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=5230 $D=1
M617 531 78 243 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=9860 $D=1
M618 247 79 529 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=600 $D=1
M619 248 79 530 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=5230 $D=1
M620 249 79 531 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=9860 $D=1
M621 532 79 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=600 $D=1
M622 533 79 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=5230 $D=1
M623 534 79 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=9860 $D=1
M624 7 80 535 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=600 $D=1
M625 7 80 536 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=5230 $D=1
M626 7 80 537 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=9860 $D=1
M627 538 81 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=600 $D=1
M628 539 81 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=5230 $D=1
M629 540 81 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=9860 $D=1
M630 541 80 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=600 $D=1
M631 542 80 227 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=5230 $D=1
M632 543 80 228 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=9860 $D=1
M633 7 541 1005 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=600 $D=1
M634 7 542 1006 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=5230 $D=1
M635 7 543 1007 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=9860 $D=1
M636 544 1005 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=600 $D=1
M637 545 1006 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=5230 $D=1
M638 546 1007 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=9860 $D=1
M639 541 535 544 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=600 $D=1
M640 542 536 545 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=5230 $D=1
M641 543 537 546 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=9860 $D=1
M642 544 81 241 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=600 $D=1
M643 545 81 242 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=5230 $D=1
M644 546 81 243 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=9860 $D=1
M645 247 82 544 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=600 $D=1
M646 248 82 545 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=5230 $D=1
M647 249 82 546 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=9860 $D=1
M648 547 82 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=600 $D=1
M649 548 82 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=5230 $D=1
M650 549 82 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=9860 $D=1
M651 7 83 550 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=600 $D=1
M652 7 83 551 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=5230 $D=1
M653 7 83 552 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=9860 $D=1
M654 553 84 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=600 $D=1
M655 554 84 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=5230 $D=1
M656 555 84 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=9860 $D=1
M657 556 83 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=600 $D=1
M658 557 83 227 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=5230 $D=1
M659 558 83 228 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=9860 $D=1
M660 7 556 1008 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=600 $D=1
M661 7 557 1009 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=5230 $D=1
M662 7 558 1010 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=9860 $D=1
M663 559 1008 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=600 $D=1
M664 560 1009 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=5230 $D=1
M665 561 1010 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=9860 $D=1
M666 556 550 559 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=600 $D=1
M667 557 551 560 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=5230 $D=1
M668 558 552 561 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=9860 $D=1
M669 559 84 241 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=600 $D=1
M670 560 84 242 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=5230 $D=1
M671 561 84 243 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=9860 $D=1
M672 247 85 559 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=600 $D=1
M673 248 85 560 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=5230 $D=1
M674 249 85 561 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=9860 $D=1
M675 562 85 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=600 $D=1
M676 563 85 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=5230 $D=1
M677 564 85 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=9860 $D=1
M678 7 86 565 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=600 $D=1
M679 7 86 566 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=5230 $D=1
M680 7 86 567 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=9860 $D=1
M681 568 87 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=600 $D=1
M682 569 87 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=5230 $D=1
M683 570 87 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=9860 $D=1
M684 571 86 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=600 $D=1
M685 572 86 227 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=5230 $D=1
M686 573 86 228 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=9860 $D=1
M687 7 571 1011 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=600 $D=1
M688 7 572 1012 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=5230 $D=1
M689 7 573 1013 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=9860 $D=1
M690 574 1011 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=600 $D=1
M691 575 1012 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=5230 $D=1
M692 576 1013 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=9860 $D=1
M693 571 565 574 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=600 $D=1
M694 572 566 575 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=5230 $D=1
M695 573 567 576 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=9860 $D=1
M696 574 87 241 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=600 $D=1
M697 575 87 242 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=5230 $D=1
M698 576 87 243 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=9860 $D=1
M699 247 88 574 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=600 $D=1
M700 248 88 575 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=5230 $D=1
M701 249 88 576 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=9860 $D=1
M702 577 88 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=600 $D=1
M703 578 88 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=5230 $D=1
M704 579 88 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=9860 $D=1
M705 7 89 580 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=600 $D=1
M706 7 89 581 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=5230 $D=1
M707 7 89 582 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=9860 $D=1
M708 583 90 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=600 $D=1
M709 584 90 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=5230 $D=1
M710 585 90 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=9860 $D=1
M711 586 89 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=600 $D=1
M712 587 89 227 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=5230 $D=1
M713 588 89 228 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=9860 $D=1
M714 7 586 1014 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=600 $D=1
M715 7 587 1015 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=5230 $D=1
M716 7 588 1016 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=9860 $D=1
M717 589 1014 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=600 $D=1
M718 590 1015 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=5230 $D=1
M719 591 1016 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=9860 $D=1
M720 586 580 589 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=600 $D=1
M721 587 581 590 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=5230 $D=1
M722 588 582 591 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=9860 $D=1
M723 589 90 241 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=600 $D=1
M724 590 90 242 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=5230 $D=1
M725 591 90 243 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=9860 $D=1
M726 247 91 589 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=600 $D=1
M727 248 91 590 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=5230 $D=1
M728 249 91 591 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=9860 $D=1
M729 592 91 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=600 $D=1
M730 593 91 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=5230 $D=1
M731 594 91 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=9860 $D=1
M732 7 92 595 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=600 $D=1
M733 7 92 596 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=5230 $D=1
M734 7 92 597 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=9860 $D=1
M735 598 93 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=600 $D=1
M736 599 93 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=5230 $D=1
M737 600 93 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=9860 $D=1
M738 601 92 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=600 $D=1
M739 602 92 227 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=5230 $D=1
M740 603 92 228 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=9860 $D=1
M741 7 601 1017 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=600 $D=1
M742 7 602 1018 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=5230 $D=1
M743 7 603 1019 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=9860 $D=1
M744 604 1017 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=600 $D=1
M745 605 1018 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=5230 $D=1
M746 606 1019 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=9860 $D=1
M747 601 595 604 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=600 $D=1
M748 602 596 605 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=5230 $D=1
M749 603 597 606 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=9860 $D=1
M750 604 93 241 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=600 $D=1
M751 605 93 242 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=5230 $D=1
M752 606 93 243 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=9860 $D=1
M753 247 94 604 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=600 $D=1
M754 248 94 605 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=5230 $D=1
M755 249 94 606 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=9860 $D=1
M756 607 94 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=600 $D=1
M757 608 94 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=5230 $D=1
M758 609 94 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=9860 $D=1
M759 7 95 610 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=600 $D=1
M760 7 95 611 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=5230 $D=1
M761 7 95 612 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=9860 $D=1
M762 613 96 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=600 $D=1
M763 614 96 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=5230 $D=1
M764 615 96 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=9860 $D=1
M765 616 95 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=600 $D=1
M766 617 95 227 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=5230 $D=1
M767 618 95 228 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=9860 $D=1
M768 7 616 1020 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=600 $D=1
M769 7 617 1021 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=5230 $D=1
M770 7 618 1022 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=9860 $D=1
M771 619 1020 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=600 $D=1
M772 620 1021 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=5230 $D=1
M773 621 1022 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=9860 $D=1
M774 616 610 619 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=600 $D=1
M775 617 611 620 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=5230 $D=1
M776 618 612 621 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=9860 $D=1
M777 619 96 241 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=600 $D=1
M778 620 96 242 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=5230 $D=1
M779 621 96 243 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=9860 $D=1
M780 247 97 619 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=600 $D=1
M781 248 97 620 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=5230 $D=1
M782 249 97 621 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=9860 $D=1
M783 622 97 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=600 $D=1
M784 623 97 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=5230 $D=1
M785 624 97 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=9860 $D=1
M786 7 98 625 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=600 $D=1
M787 7 98 626 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=5230 $D=1
M788 7 98 627 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=9860 $D=1
M789 628 99 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=600 $D=1
M790 629 99 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=5230 $D=1
M791 630 99 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=9860 $D=1
M792 631 98 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=600 $D=1
M793 632 98 227 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=5230 $D=1
M794 633 98 228 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=9860 $D=1
M795 7 631 1023 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=600 $D=1
M796 7 632 1024 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=5230 $D=1
M797 7 633 1025 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=9860 $D=1
M798 634 1023 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=600 $D=1
M799 635 1024 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=5230 $D=1
M800 636 1025 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=9860 $D=1
M801 631 625 634 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=600 $D=1
M802 632 626 635 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=5230 $D=1
M803 633 627 636 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=9860 $D=1
M804 634 99 241 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=600 $D=1
M805 635 99 242 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=5230 $D=1
M806 636 99 243 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=9860 $D=1
M807 247 100 634 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=600 $D=1
M808 248 100 635 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=5230 $D=1
M809 249 100 636 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=9860 $D=1
M810 637 100 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=600 $D=1
M811 638 100 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=5230 $D=1
M812 639 100 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=9860 $D=1
M813 7 101 640 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=600 $D=1
M814 7 101 641 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=5230 $D=1
M815 7 101 642 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=9860 $D=1
M816 643 102 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=600 $D=1
M817 644 102 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=5230 $D=1
M818 645 102 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=9860 $D=1
M819 646 101 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=600 $D=1
M820 647 101 227 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=5230 $D=1
M821 648 101 228 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=9860 $D=1
M822 7 646 1026 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=600 $D=1
M823 7 647 1027 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=5230 $D=1
M824 7 648 1028 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=9860 $D=1
M825 649 1026 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=600 $D=1
M826 650 1027 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=5230 $D=1
M827 651 1028 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=9860 $D=1
M828 646 640 649 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=600 $D=1
M829 647 641 650 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=5230 $D=1
M830 648 642 651 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=9860 $D=1
M831 649 102 241 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=600 $D=1
M832 650 102 242 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=5230 $D=1
M833 651 102 243 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=9860 $D=1
M834 247 103 649 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=600 $D=1
M835 248 103 650 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=5230 $D=1
M836 249 103 651 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=9860 $D=1
M837 652 103 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=600 $D=1
M838 653 103 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=5230 $D=1
M839 654 103 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=9860 $D=1
M840 7 104 655 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=600 $D=1
M841 7 104 656 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=5230 $D=1
M842 7 104 657 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=9860 $D=1
M843 658 105 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=600 $D=1
M844 659 105 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=5230 $D=1
M845 660 105 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=9860 $D=1
M846 661 104 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=600 $D=1
M847 662 104 227 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=5230 $D=1
M848 663 104 228 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=9860 $D=1
M849 7 661 1029 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=600 $D=1
M850 7 662 1030 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=5230 $D=1
M851 7 663 1031 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=9860 $D=1
M852 664 1029 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=600 $D=1
M853 665 1030 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=5230 $D=1
M854 666 1031 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=9860 $D=1
M855 661 655 664 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=600 $D=1
M856 662 656 665 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=5230 $D=1
M857 663 657 666 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=9860 $D=1
M858 664 105 241 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=600 $D=1
M859 665 105 242 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=5230 $D=1
M860 666 105 243 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=9860 $D=1
M861 247 106 664 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=600 $D=1
M862 248 106 665 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=5230 $D=1
M863 249 106 666 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=9860 $D=1
M864 667 106 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=600 $D=1
M865 668 106 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=5230 $D=1
M866 669 106 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=9860 $D=1
M867 7 107 670 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=600 $D=1
M868 7 107 671 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=5230 $D=1
M869 7 107 672 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=9860 $D=1
M870 673 108 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=600 $D=1
M871 674 108 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=5230 $D=1
M872 675 108 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=9860 $D=1
M873 676 107 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=600 $D=1
M874 677 107 227 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=5230 $D=1
M875 678 107 228 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=9860 $D=1
M876 7 676 1032 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=600 $D=1
M877 7 677 1033 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=5230 $D=1
M878 7 678 1034 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=9860 $D=1
M879 679 1032 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=600 $D=1
M880 680 1033 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=5230 $D=1
M881 681 1034 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=9860 $D=1
M882 676 670 679 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=600 $D=1
M883 677 671 680 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=5230 $D=1
M884 678 672 681 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=9860 $D=1
M885 679 108 241 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=600 $D=1
M886 680 108 242 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=5230 $D=1
M887 681 108 243 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=9860 $D=1
M888 247 111 679 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=600 $D=1
M889 248 111 680 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=5230 $D=1
M890 249 111 681 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=9860 $D=1
M891 682 111 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=600 $D=1
M892 683 111 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=5230 $D=1
M893 684 111 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=9860 $D=1
M894 7 112 685 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=600 $D=1
M895 7 112 686 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=5230 $D=1
M896 7 112 687 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=9860 $D=1
M897 688 113 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=600 $D=1
M898 689 113 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=5230 $D=1
M899 690 113 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=9860 $D=1
M900 691 112 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=600 $D=1
M901 692 112 227 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=5230 $D=1
M902 693 112 228 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=9860 $D=1
M903 7 691 1035 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=600 $D=1
M904 7 692 1036 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=5230 $D=1
M905 7 693 1037 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=9860 $D=1
M906 694 1035 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=600 $D=1
M907 695 1036 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=5230 $D=1
M908 696 1037 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=9860 $D=1
M909 691 685 694 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=600 $D=1
M910 692 686 695 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=5230 $D=1
M911 693 687 696 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=9860 $D=1
M912 694 113 241 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=600 $D=1
M913 695 113 242 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=5230 $D=1
M914 696 113 243 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=9860 $D=1
M915 247 116 694 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=600 $D=1
M916 248 116 695 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=5230 $D=1
M917 249 116 696 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=9860 $D=1
M918 697 116 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=600 $D=1
M919 698 116 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=5230 $D=1
M920 699 116 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=9860 $D=1
M921 7 117 700 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=600 $D=1
M922 7 117 701 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=5230 $D=1
M923 7 117 702 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=9860 $D=1
M924 703 118 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=600 $D=1
M925 704 118 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=5230 $D=1
M926 705 118 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=9860 $D=1
M927 7 118 241 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=600 $D=1
M928 7 118 242 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=5230 $D=1
M929 7 118 243 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=9860 $D=1
M930 247 117 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=600 $D=1
M931 248 117 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=5230 $D=1
M932 249 117 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=9860 $D=1
M933 7 709 706 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=600 $D=1
M934 7 710 707 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=5230 $D=1
M935 7 711 708 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=9860 $D=1
M936 709 119 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=600 $D=1
M937 710 119 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=5230 $D=1
M938 711 119 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=9860 $D=1
M939 1038 241 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=600 $D=1
M940 1039 242 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=5230 $D=1
M941 1040 243 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=9860 $D=1
M942 712 706 1038 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=600 $D=1
M943 713 707 1039 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=5230 $D=1
M944 714 708 1040 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=9860 $D=1
M945 7 712 120 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=600 $D=1
M946 7 713 715 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=5230 $D=1
M947 7 714 716 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=9860 $D=1
M948 1041 120 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=600 $D=1
M949 1042 715 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=5230 $D=1
M950 1043 716 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=9860 $D=1
M951 712 709 1041 7 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=600 $D=1
M952 713 710 1042 7 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=5230 $D=1
M953 714 711 1043 7 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=9860 $D=1
M954 7 720 717 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=600 $D=1
M955 7 721 718 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=5230 $D=1
M956 7 722 719 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=9860 $D=1
M957 720 119 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=600 $D=1
M958 721 119 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=5230 $D=1
M959 722 119 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=9860 $D=1
M960 1044 247 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=600 $D=1
M961 1045 248 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=5230 $D=1
M962 1046 249 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=9860 $D=1
M963 723 717 1044 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=600 $D=1
M964 724 718 1045 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=5230 $D=1
M965 725 719 1046 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=9860 $D=1
M966 7 723 121 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=600 $D=1
M967 7 724 122 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=5230 $D=1
M968 7 725 123 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=9860 $D=1
M969 1047 121 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=600 $D=1
M970 1048 122 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=5230 $D=1
M971 1049 123 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=9860 $D=1
M972 723 720 1047 7 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=600 $D=1
M973 724 721 1048 7 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=5230 $D=1
M974 725 722 1049 7 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=9860 $D=1
M975 726 124 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=600 $D=1
M976 727 124 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=5230 $D=1
M977 728 124 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=9860 $D=1
M978 729 726 120 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=600 $D=1
M979 730 727 715 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=5230 $D=1
M980 731 728 716 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=9860 $D=1
M981 125 124 729 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=600 $D=1
M982 126 124 730 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=5230 $D=1
M983 127 124 731 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=9860 $D=1
M984 732 128 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=600 $D=1
M985 733 128 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=5230 $D=1
M986 734 128 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=9860 $D=1
M987 735 732 121 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=600 $D=1
M988 736 733 122 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=5230 $D=1
M989 737 734 123 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=9860 $D=1
M990 1050 128 735 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=600 $D=1
M991 1051 128 736 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=5230 $D=1
M992 1052 128 737 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=9860 $D=1
M993 7 121 1050 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=600 $D=1
M994 7 122 1051 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=5230 $D=1
M995 7 123 1052 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=9860 $D=1
M996 738 129 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=600 $D=1
M997 739 129 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=5230 $D=1
M998 740 129 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=9860 $D=1
M999 741 738 735 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=600 $D=1
M1000 742 739 736 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=5230 $D=1
M1001 743 740 737 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=9860 $D=1
M1002 12 129 741 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=600 $D=1
M1003 13 129 742 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=5230 $D=1
M1004 14 129 743 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=9860 $D=1
M1005 746 744 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=600 $D=1
M1006 747 745 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=5230 $D=1
M1007 748 130 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=9860 $D=1
M1008 7 752 749 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=600 $D=1
M1009 7 753 750 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=5230 $D=1
M1010 7 754 751 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=9860 $D=1
M1011 755 729 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=600 $D=1
M1012 756 730 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=5230 $D=1
M1013 757 731 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=9860 $D=1
M1014 752 755 744 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=600 $D=1
M1015 753 756 745 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=5230 $D=1
M1016 754 757 130 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=9860 $D=1
M1017 746 729 752 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=600 $D=1
M1018 747 730 753 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=5230 $D=1
M1019 748 731 754 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=9860 $D=1
M1020 758 749 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=600 $D=1
M1021 759 750 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=5230 $D=1
M1022 760 751 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=9860 $D=1
M1023 761 758 741 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=600 $D=1
M1024 744 759 742 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=5230 $D=1
M1025 745 760 743 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=9860 $D=1
M1026 729 749 761 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=600 $D=1
M1027 730 750 744 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=5230 $D=1
M1028 731 751 745 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=9860 $D=1
M1029 762 761 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=600 $D=1
M1030 763 744 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=5230 $D=1
M1031 764 745 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=9860 $D=1
M1032 765 749 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=600 $D=1
M1033 766 750 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=5230 $D=1
M1034 767 751 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=9860 $D=1
M1035 768 765 762 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=600 $D=1
M1036 769 766 763 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=5230 $D=1
M1037 770 767 764 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=9860 $D=1
M1038 741 749 768 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=600 $D=1
M1039 742 750 769 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=5230 $D=1
M1040 743 751 770 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=9860 $D=1
M1041 771 729 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=600 $D=1
M1042 772 730 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=5230 $D=1
M1043 773 731 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=9860 $D=1
M1044 7 741 771 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=600 $D=1
M1045 7 742 772 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=5230 $D=1
M1046 7 743 773 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=9860 $D=1
M1047 774 768 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=600 $D=1
M1048 775 769 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=5230 $D=1
M1049 776 770 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=9860 $D=1
M1050 1080 729 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=600 $D=1
M1051 1081 730 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=5230 $D=1
M1052 1082 731 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=9860 $D=1
M1053 777 741 1080 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=600 $D=1
M1054 778 742 1081 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=5230 $D=1
M1055 779 743 1082 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=9860 $D=1
M1056 1083 729 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=600 $D=1
M1057 1084 730 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=5230 $D=1
M1058 1085 731 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=9860 $D=1
M1059 780 741 1083 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=600 $D=1
M1060 781 742 1084 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=5230 $D=1
M1061 782 743 1085 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=9860 $D=1
M1062 786 729 783 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=600 $D=1
M1063 787 730 784 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=5230 $D=1
M1064 788 731 785 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=9860 $D=1
M1065 783 741 786 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=600 $D=1
M1066 784 742 787 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=5230 $D=1
M1067 785 743 788 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=9860 $D=1
M1068 7 780 783 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=600 $D=1
M1069 7 781 784 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=5230 $D=1
M1070 7 782 785 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=9860 $D=1
M1071 789 134 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=600 $D=1
M1072 790 134 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=5230 $D=1
M1073 791 134 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=9860 $D=1
M1074 792 789 771 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=600 $D=1
M1075 793 790 772 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=5230 $D=1
M1076 794 791 773 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=9860 $D=1
M1077 777 134 792 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=600 $D=1
M1078 778 134 793 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=5230 $D=1
M1079 779 134 794 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=9860 $D=1
M1080 795 789 774 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=600 $D=1
M1081 796 790 775 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=5230 $D=1
M1082 797 791 776 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=9860 $D=1
M1083 786 134 795 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=600 $D=1
M1084 787 134 796 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=5230 $D=1
M1085 788 134 797 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=9860 $D=1
M1086 798 135 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=600 $D=1
M1087 799 135 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=5230 $D=1
M1088 800 135 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=9860 $D=1
M1089 801 798 795 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=600 $D=1
M1090 802 799 796 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=5230 $D=1
M1091 803 800 797 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=9860 $D=1
M1092 792 135 801 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=600 $D=1
M1093 793 135 802 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=5230 $D=1
M1094 794 135 803 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=9860 $D=1
M1095 15 801 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=600 $D=1
M1096 16 802 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=5230 $D=1
M1097 17 803 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=9860 $D=1
M1098 804 136 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=600 $D=1
M1099 805 136 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=5230 $D=1
M1100 806 136 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=9860 $D=1
M1101 808 804 807 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=600 $D=1
M1102 809 805 137 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=5230 $D=1
M1103 810 806 138 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=9860 $D=1
M1104 139 136 808 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=600 $D=1
M1105 811 136 809 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=5230 $D=1
M1106 807 136 810 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=9860 $D=1
M1107 812 136 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=600 $D=1
M1108 813 136 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=5230 $D=1
M1109 814 136 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=9860 $D=1
M1110 815 812 140 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=600 $D=1
M1111 816 813 141 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=5230 $D=1
M1112 817 814 142 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=9860 $D=1
M1113 139 136 815 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=600 $D=1
M1114 139 136 816 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=5230 $D=1
M1115 818 136 817 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=9860 $D=1
M1116 819 136 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=600 $D=1
M1117 820 136 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=5230 $D=1
M1118 821 136 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=9860 $D=1
M1119 822 819 133 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=600 $D=1
M1120 823 820 132 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=5230 $D=1
M1121 824 821 131 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=9860 $D=1
M1122 139 136 822 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=600 $D=1
M1123 139 136 823 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=5230 $D=1
M1124 139 136 824 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=9860 $D=1
M1125 825 136 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=600 $D=1
M1126 826 136 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=5230 $D=1
M1127 827 136 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=9860 $D=1
M1128 828 825 143 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=600 $D=1
M1129 829 826 144 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=5230 $D=1
M1130 830 827 145 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=9860 $D=1
M1131 139 136 828 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=600 $D=1
M1132 139 136 829 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=5230 $D=1
M1133 139 136 830 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=9860 $D=1
M1134 831 136 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=600 $D=1
M1135 832 136 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=5230 $D=1
M1136 833 136 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=9860 $D=1
M1137 834 831 146 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=600 $D=1
M1138 835 832 147 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=5230 $D=1
M1139 836 833 148 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=9860 $D=1
M1140 139 136 834 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=600 $D=1
M1141 139 136 835 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=5230 $D=1
M1142 139 136 836 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=9860 $D=1
M1143 7 729 1053 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=600 $D=1
M1144 7 730 1054 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=5230 $D=1
M1145 7 731 1055 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=9860 $D=1
M1146 811 1053 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=600 $D=1
M1147 807 1054 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=5230 $D=1
M1148 137 1055 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=9860 $D=1
M1149 837 149 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=600 $D=1
M1150 838 149 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=5230 $D=1
M1151 839 149 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=9860 $D=1
M1152 818 837 811 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=600 $D=1
M1153 150 838 807 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=5230 $D=1
M1154 140 839 137 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=9860 $D=1
M1155 808 149 818 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=600 $D=1
M1156 809 149 150 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=5230 $D=1
M1157 810 149 140 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=9860 $D=1
M1158 840 151 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=600 $D=1
M1159 841 151 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=5230 $D=1
M1160 842 151 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=9860 $D=1
M1161 152 840 818 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=600 $D=1
M1162 153 841 150 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=5230 $D=1
M1163 154 842 140 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=9860 $D=1
M1164 815 151 152 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=600 $D=1
M1165 816 151 153 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=5230 $D=1
M1166 817 151 154 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=9860 $D=1
M1167 843 155 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=600 $D=1
M1168 844 155 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=5230 $D=1
M1169 845 155 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=9860 $D=1
M1170 110 843 152 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=600 $D=1
M1171 114 844 153 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=5230 $D=1
M1172 109 845 154 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=9860 $D=1
M1173 822 155 110 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=600 $D=1
M1174 823 155 114 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=5230 $D=1
M1175 824 155 109 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=9860 $D=1
M1176 846 156 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=600 $D=1
M1177 847 156 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=5230 $D=1
M1178 848 156 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=9860 $D=1
M1179 157 846 110 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=600 $D=1
M1180 158 847 114 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=5230 $D=1
M1181 159 848 109 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=9860 $D=1
M1182 828 156 157 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=600 $D=1
M1183 829 156 158 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=5230 $D=1
M1184 830 156 159 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=9860 $D=1
M1185 849 160 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=600 $D=1
M1186 850 160 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=5230 $D=1
M1187 851 160 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=9860 $D=1
M1188 205 849 157 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=600 $D=1
M1189 206 850 158 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=5230 $D=1
M1190 207 851 159 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=9860 $D=1
M1191 834 160 205 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=600 $D=1
M1192 835 160 206 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=5230 $D=1
M1193 836 160 207 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=9860 $D=1
M1194 852 161 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=600 $D=1
M1195 853 161 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=5230 $D=1
M1196 854 161 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=9860 $D=1
M1197 162 852 121 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=600 $D=1
M1198 855 853 122 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=5230 $D=1
M1199 856 854 123 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=9860 $D=1
M1200 12 161 162 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=600 $D=1
M1201 13 161 855 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=5230 $D=1
M1202 14 161 856 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=9860 $D=1
M1203 1086 120 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=600 $D=1
M1204 1087 715 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=5230 $D=1
M1205 1088 716 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=9860 $D=1
M1206 857 162 1086 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=600 $D=1
M1207 858 855 1087 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=5230 $D=1
M1208 859 856 1088 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=9860 $D=1
M1209 863 120 860 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=600 $D=1
M1210 864 715 861 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=5230 $D=1
M1211 865 716 862 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=9860 $D=1
M1212 860 162 863 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=600 $D=1
M1213 861 855 864 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=5230 $D=1
M1214 862 856 865 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=9860 $D=1
M1215 7 857 860 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=600 $D=1
M1216 7 858 861 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=5230 $D=1
M1217 7 859 862 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=9860 $D=1
M1218 1089 10 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=600 $D=1
M1219 1090 866 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=5230 $D=1
M1220 1091 867 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=9860 $D=1
M1221 1056 863 1089 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=600 $D=1
M1222 1057 864 1090 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=5230 $D=1
M1223 1058 865 1091 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=9860 $D=1
M1224 866 1056 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=600 $D=1
M1225 867 1057 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=5230 $D=1
M1226 163 1058 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=9860 $D=1
M1227 868 120 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=600 $D=1
M1228 869 715 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=5230 $D=1
M1229 870 716 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=9860 $D=1
M1230 7 871 868 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=600 $D=1
M1231 7 872 869 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=5230 $D=1
M1232 7 873 870 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=9860 $D=1
M1233 871 162 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=600 $D=1
M1234 872 855 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=5230 $D=1
M1235 873 856 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=9860 $D=1
M1236 1092 868 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=600 $D=1
M1237 1093 869 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=5230 $D=1
M1238 1094 870 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=9860 $D=1
M1239 874 10 1092 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=600 $D=1
M1240 875 866 1093 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=5230 $D=1
M1241 876 867 1094 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=9860 $D=1
M1242 879 7 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=600 $D=1
M1243 880 877 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=5230 $D=1
M1244 881 878 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=9860 $D=1
M1245 1095 874 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=600 $D=1
M1246 1096 875 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=5230 $D=1
M1247 1097 876 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=9860 $D=1
M1248 877 879 1095 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=600 $D=1
M1249 878 880 1096 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=5230 $D=1
M1250 164 881 1097 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=9860 $D=1
M1251 884 882 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=600 $D=1
M1252 885 883 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=5230 $D=1
M1253 886 165 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=9860 $D=1
M1254 7 890 887 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=600 $D=1
M1255 7 891 888 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=5230 $D=1
M1256 7 892 889 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=9860 $D=1
M1257 893 125 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=600 $D=1
M1258 894 126 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=5230 $D=1
M1259 895 127 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=9860 $D=1
M1260 890 893 882 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=600 $D=1
M1261 891 894 883 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=5230 $D=1
M1262 892 895 165 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=9860 $D=1
M1263 884 125 890 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=600 $D=1
M1264 885 126 891 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=5230 $D=1
M1265 886 127 892 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=9860 $D=1
M1266 896 887 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=600 $D=1
M1267 897 888 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=5230 $D=1
M1268 898 889 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=9860 $D=1
M1269 899 896 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=600 $D=1
M1270 882 897 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=5230 $D=1
M1271 883 898 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=9860 $D=1
M1272 125 887 899 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=600 $D=1
M1273 126 888 882 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=5230 $D=1
M1274 127 889 883 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=9860 $D=1
M1275 900 899 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=600 $D=1
M1276 901 882 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=5230 $D=1
M1277 902 883 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=9860 $D=1
M1278 903 887 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=600 $D=1
M1279 904 888 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=5230 $D=1
M1280 905 889 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=9860 $D=1
M1281 208 903 900 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=600 $D=1
M1282 209 904 901 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=5230 $D=1
M1283 210 905 902 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=9860 $D=1
M1284 7 887 208 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=600 $D=1
M1285 7 888 209 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=5230 $D=1
M1286 7 889 210 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=9860 $D=1
M1287 906 166 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=600 $D=1
M1288 907 166 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=5230 $D=1
M1289 908 166 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=9860 $D=1
M1290 909 906 208 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=600 $D=1
M1291 910 907 209 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=5230 $D=1
M1292 911 908 210 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=9860 $D=1
M1293 15 166 909 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=600 $D=1
M1294 16 166 910 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=5230 $D=1
M1295 17 166 911 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=9860 $D=1
M1296 912 167 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=600 $D=1
M1297 913 167 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=5230 $D=1
M1298 914 167 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=9860 $D=1
M1299 915 912 909 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=600 $D=1
M1300 916 913 910 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=5230 $D=1
M1301 917 914 911 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=9860 $D=1
M1302 7 167 915 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=600 $D=1
M1303 10 167 916 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=5230 $D=1
M1304 10 167 917 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=9860 $D=1
M1305 918 119 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=600 $D=1
M1306 919 119 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=5230 $D=1
M1307 920 119 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=9860 $D=1
M1308 7 918 921 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=600 $D=1
M1309 7 919 922 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=5230 $D=1
M1310 7 920 923 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=9860 $D=1
M1311 924 119 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=600 $D=1
M1312 925 119 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=5230 $D=1
M1313 926 119 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=9860 $D=1
M1314 927 918 915 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=600 $D=1
M1315 928 919 916 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=5230 $D=1
M1316 929 920 917 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=9860 $D=1
M1317 7 927 1059 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=600 $D=1
M1318 7 928 1060 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=5230 $D=1
M1319 7 929 1061 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=9860 $D=1
M1320 930 1059 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=600 $D=1
M1321 931 1060 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=5230 $D=1
M1322 932 1061 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=9860 $D=1
M1323 927 921 930 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=600 $D=1
M1324 928 922 931 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=5230 $D=1
M1325 929 923 932 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=9860 $D=1
M1326 933 119 930 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=600 $D=1
M1327 934 119 931 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=5230 $D=1
M1328 935 119 932 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=9860 $D=1
M1329 7 939 936 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=600 $D=1
M1330 7 940 937 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=5230 $D=1
M1331 7 941 938 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=9860 $D=1
M1332 939 119 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=600 $D=1
M1333 940 119 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=5230 $D=1
M1334 941 119 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=9860 $D=1
M1335 1062 933 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=600 $D=1
M1336 1063 934 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=5230 $D=1
M1337 1064 935 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=9860 $D=1
M1338 942 936 1062 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=600 $D=1
M1339 943 937 1063 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=5230 $D=1
M1340 944 938 1064 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=9860 $D=1
M1341 7 942 125 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=600 $D=1
M1342 7 943 126 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=5230 $D=1
M1343 7 944 127 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=9860 $D=1
M1344 1065 125 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=600 $D=1
M1345 1066 126 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=5230 $D=1
M1346 1067 127 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=9860 $D=1
M1347 942 939 1065 7 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=600 $D=1
M1348 943 940 1066 7 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=5230 $D=1
M1349 944 941 1067 7 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=9860 $D=1
M1350 169 1 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=1850 $D=0
M1351 170 1 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=6480 $D=0
M1352 171 1 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=11110 $D=0
M1353 172 1 2 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=1850 $D=0
M1354 173 1 3 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=6480 $D=0
M1355 174 1 4 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=11110 $D=0
M1356 7 169 172 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=1850 $D=0
M1357 7 170 173 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=6480 $D=0
M1358 7 171 174 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=11110 $D=0
M1359 175 1 5 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=1850 $D=0
M1360 176 1 5 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=6480 $D=0
M1361 177 1 5 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=11110 $D=0
M1362 6 169 175 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=1850 $D=0
M1363 6 170 176 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=6480 $D=0
M1364 6 171 177 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=11110 $D=0
M1365 178 1 7 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=1850 $D=0
M1366 179 1 7 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=6480 $D=0
M1367 180 1 7 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=11110 $D=0
M1368 7 169 178 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=1850 $D=0
M1369 7 170 179 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=6480 $D=0
M1370 7 171 180 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=11110 $D=0
M1371 184 8 178 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=1850 $D=0
M1372 185 8 179 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=6480 $D=0
M1373 186 8 180 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=11110 $D=0
M1374 181 8 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=1850 $D=0
M1375 182 8 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=6480 $D=0
M1376 183 8 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=11110 $D=0
M1377 187 8 175 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=1850 $D=0
M1378 188 8 176 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=6480 $D=0
M1379 189 8 177 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=11110 $D=0
M1380 172 181 187 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=1850 $D=0
M1381 173 182 188 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=6480 $D=0
M1382 174 183 189 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=11110 $D=0
M1383 190 9 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=1850 $D=0
M1384 191 9 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=6480 $D=0
M1385 192 9 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=11110 $D=0
M1386 193 9 187 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=1850 $D=0
M1387 194 9 188 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=6480 $D=0
M1388 195 9 189 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=11110 $D=0
M1389 184 190 193 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=1850 $D=0
M1390 185 191 194 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=6480 $D=0
M1391 186 192 195 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=11110 $D=0
M1392 196 11 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=1850 $D=0
M1393 197 11 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=6480 $D=0
M1394 198 11 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=11110 $D=0
M1395 199 11 7 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=1850 $D=0
M1396 200 11 7 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=6480 $D=0
M1397 201 11 7 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=11110 $D=0
M1398 12 196 199 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=1850 $D=0
M1399 13 197 200 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=6480 $D=0
M1400 14 198 201 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=11110 $D=0
M1401 202 11 15 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=1850 $D=0
M1402 203 11 16 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=6480 $D=0
M1403 204 11 17 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=11110 $D=0
M1404 205 196 202 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=1850 $D=0
M1405 206 197 203 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=6480 $D=0
M1406 207 198 204 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=11110 $D=0
M1407 211 11 208 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=1850 $D=0
M1408 212 11 209 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=6480 $D=0
M1409 213 11 210 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=11110 $D=0
M1410 193 196 211 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=1850 $D=0
M1411 194 197 212 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=6480 $D=0
M1412 195 198 213 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=11110 $D=0
M1413 217 18 211 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=1850 $D=0
M1414 218 18 212 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=6480 $D=0
M1415 219 18 213 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=11110 $D=0
M1416 214 18 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=1850 $D=0
M1417 215 18 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=6480 $D=0
M1418 216 18 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=11110 $D=0
M1419 220 18 202 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=1850 $D=0
M1420 221 18 203 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=6480 $D=0
M1421 222 18 204 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=11110 $D=0
M1422 199 214 220 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=1850 $D=0
M1423 200 215 221 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=6480 $D=0
M1424 201 216 222 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=11110 $D=0
M1425 223 19 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=1850 $D=0
M1426 224 19 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=6480 $D=0
M1427 225 19 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=11110 $D=0
M1428 226 19 220 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=1850 $D=0
M1429 227 19 221 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=6480 $D=0
M1430 228 19 222 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=11110 $D=0
M1431 217 223 226 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=1850 $D=0
M1432 218 224 227 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=6480 $D=0
M1433 219 225 228 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=11110 $D=0
M1434 10 20 229 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=1850 $D=0
M1435 10 20 230 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=6480 $D=0
M1436 10 20 231 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=11110 $D=0
M1437 232 21 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=1850 $D=0
M1438 233 21 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=6480 $D=0
M1439 234 21 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=11110 $D=0
M1440 235 229 226 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=1850 $D=0
M1441 236 230 227 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=6480 $D=0
M1442 237 231 228 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=11110 $D=0
M1443 10 235 945 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=1850 $D=0
M1444 10 236 946 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=6480 $D=0
M1445 10 237 947 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=11110 $D=0
M1446 238 945 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=1850 $D=0
M1447 239 946 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=6480 $D=0
M1448 240 947 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=11110 $D=0
M1449 235 20 238 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=1850 $D=0
M1450 236 20 239 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=6480 $D=0
M1451 237 20 240 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=11110 $D=0
M1452 238 232 241 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=1850 $D=0
M1453 239 233 242 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=6480 $D=0
M1454 240 234 243 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=11110 $D=0
M1455 247 244 238 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=1850 $D=0
M1456 248 245 239 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=6480 $D=0
M1457 249 246 240 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=11110 $D=0
M1458 244 22 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=1850 $D=0
M1459 245 22 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=6480 $D=0
M1460 246 22 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=11110 $D=0
M1461 10 23 250 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=1850 $D=0
M1462 10 23 251 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=6480 $D=0
M1463 10 23 252 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=11110 $D=0
M1464 253 24 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=1850 $D=0
M1465 254 24 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=6480 $D=0
M1466 255 24 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=11110 $D=0
M1467 256 250 226 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=1850 $D=0
M1468 257 251 227 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=6480 $D=0
M1469 258 252 228 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=11110 $D=0
M1470 10 256 948 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=1850 $D=0
M1471 10 257 949 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=6480 $D=0
M1472 10 258 950 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=11110 $D=0
M1473 259 948 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=1850 $D=0
M1474 260 949 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=6480 $D=0
M1475 261 950 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=11110 $D=0
M1476 256 23 259 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=1850 $D=0
M1477 257 23 260 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=6480 $D=0
M1478 258 23 261 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=11110 $D=0
M1479 259 253 241 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=1850 $D=0
M1480 260 254 242 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=6480 $D=0
M1481 261 255 243 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=11110 $D=0
M1482 247 262 259 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=1850 $D=0
M1483 248 263 260 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=6480 $D=0
M1484 249 264 261 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=11110 $D=0
M1485 262 25 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=1850 $D=0
M1486 263 25 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=6480 $D=0
M1487 264 25 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=11110 $D=0
M1488 10 26 265 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=1850 $D=0
M1489 10 26 266 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=6480 $D=0
M1490 10 26 267 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=11110 $D=0
M1491 268 27 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=1850 $D=0
M1492 269 27 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=6480 $D=0
M1493 270 27 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=11110 $D=0
M1494 271 265 226 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=1850 $D=0
M1495 272 266 227 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=6480 $D=0
M1496 273 267 228 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=11110 $D=0
M1497 10 271 951 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=1850 $D=0
M1498 10 272 952 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=6480 $D=0
M1499 10 273 953 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=11110 $D=0
M1500 274 951 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=1850 $D=0
M1501 275 952 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=6480 $D=0
M1502 276 953 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=11110 $D=0
M1503 271 26 274 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=1850 $D=0
M1504 272 26 275 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=6480 $D=0
M1505 273 26 276 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=11110 $D=0
M1506 274 268 241 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=1850 $D=0
M1507 275 269 242 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=6480 $D=0
M1508 276 270 243 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=11110 $D=0
M1509 247 277 274 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=1850 $D=0
M1510 248 278 275 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=6480 $D=0
M1511 249 279 276 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=11110 $D=0
M1512 277 28 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=1850 $D=0
M1513 278 28 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=6480 $D=0
M1514 279 28 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=11110 $D=0
M1515 10 29 280 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=1850 $D=0
M1516 10 29 281 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=6480 $D=0
M1517 10 29 282 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=11110 $D=0
M1518 283 30 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=1850 $D=0
M1519 284 30 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=6480 $D=0
M1520 285 30 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=11110 $D=0
M1521 286 280 226 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=1850 $D=0
M1522 287 281 227 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=6480 $D=0
M1523 288 282 228 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=11110 $D=0
M1524 10 286 954 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=1850 $D=0
M1525 10 287 955 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=6480 $D=0
M1526 10 288 956 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=11110 $D=0
M1527 289 954 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=1850 $D=0
M1528 290 955 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=6480 $D=0
M1529 291 956 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=11110 $D=0
M1530 286 29 289 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=1850 $D=0
M1531 287 29 290 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=6480 $D=0
M1532 288 29 291 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=11110 $D=0
M1533 289 283 241 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=1850 $D=0
M1534 290 284 242 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=6480 $D=0
M1535 291 285 243 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=11110 $D=0
M1536 247 292 289 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=1850 $D=0
M1537 248 293 290 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=6480 $D=0
M1538 249 294 291 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=11110 $D=0
M1539 292 31 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=1850 $D=0
M1540 293 31 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=6480 $D=0
M1541 294 31 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=11110 $D=0
M1542 10 32 295 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=1850 $D=0
M1543 10 32 296 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=6480 $D=0
M1544 10 32 297 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=11110 $D=0
M1545 298 33 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=1850 $D=0
M1546 299 33 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=6480 $D=0
M1547 300 33 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=11110 $D=0
M1548 301 295 226 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=1850 $D=0
M1549 302 296 227 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=6480 $D=0
M1550 303 297 228 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=11110 $D=0
M1551 10 301 957 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=1850 $D=0
M1552 10 302 958 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=6480 $D=0
M1553 10 303 959 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=11110 $D=0
M1554 304 957 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=1850 $D=0
M1555 305 958 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=6480 $D=0
M1556 306 959 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=11110 $D=0
M1557 301 32 304 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=1850 $D=0
M1558 302 32 305 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=6480 $D=0
M1559 303 32 306 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=11110 $D=0
M1560 304 298 241 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=1850 $D=0
M1561 305 299 242 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=6480 $D=0
M1562 306 300 243 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=11110 $D=0
M1563 247 307 304 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=1850 $D=0
M1564 248 308 305 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=6480 $D=0
M1565 249 309 306 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=11110 $D=0
M1566 307 34 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=1850 $D=0
M1567 308 34 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=6480 $D=0
M1568 309 34 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=11110 $D=0
M1569 10 35 310 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=1850 $D=0
M1570 10 35 311 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=6480 $D=0
M1571 10 35 312 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=11110 $D=0
M1572 313 36 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=1850 $D=0
M1573 314 36 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=6480 $D=0
M1574 315 36 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=11110 $D=0
M1575 316 310 226 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=1850 $D=0
M1576 317 311 227 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=6480 $D=0
M1577 318 312 228 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=11110 $D=0
M1578 10 316 960 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=1850 $D=0
M1579 10 317 961 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=6480 $D=0
M1580 10 318 962 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=11110 $D=0
M1581 319 960 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=1850 $D=0
M1582 320 961 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=6480 $D=0
M1583 321 962 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=11110 $D=0
M1584 316 35 319 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=1850 $D=0
M1585 317 35 320 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=6480 $D=0
M1586 318 35 321 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=11110 $D=0
M1587 319 313 241 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=1850 $D=0
M1588 320 314 242 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=6480 $D=0
M1589 321 315 243 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=11110 $D=0
M1590 247 322 319 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=1850 $D=0
M1591 248 323 320 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=6480 $D=0
M1592 249 324 321 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=11110 $D=0
M1593 322 37 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=1850 $D=0
M1594 323 37 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=6480 $D=0
M1595 324 37 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=11110 $D=0
M1596 10 38 325 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=1850 $D=0
M1597 10 38 326 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=6480 $D=0
M1598 10 38 327 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=11110 $D=0
M1599 328 39 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=1850 $D=0
M1600 329 39 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=6480 $D=0
M1601 330 39 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=11110 $D=0
M1602 331 325 226 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=1850 $D=0
M1603 332 326 227 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=6480 $D=0
M1604 333 327 228 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=11110 $D=0
M1605 10 331 963 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=1850 $D=0
M1606 10 332 964 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=6480 $D=0
M1607 10 333 965 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=11110 $D=0
M1608 334 963 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=1850 $D=0
M1609 335 964 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=6480 $D=0
M1610 336 965 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=11110 $D=0
M1611 331 38 334 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=1850 $D=0
M1612 332 38 335 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=6480 $D=0
M1613 333 38 336 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=11110 $D=0
M1614 334 328 241 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=1850 $D=0
M1615 335 329 242 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=6480 $D=0
M1616 336 330 243 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=11110 $D=0
M1617 247 337 334 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=1850 $D=0
M1618 248 338 335 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=6480 $D=0
M1619 249 339 336 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=11110 $D=0
M1620 337 40 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=1850 $D=0
M1621 338 40 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=6480 $D=0
M1622 339 40 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=11110 $D=0
M1623 10 41 340 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=1850 $D=0
M1624 10 41 341 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=6480 $D=0
M1625 10 41 342 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=11110 $D=0
M1626 343 42 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=1850 $D=0
M1627 344 42 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=6480 $D=0
M1628 345 42 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=11110 $D=0
M1629 346 340 226 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=1850 $D=0
M1630 347 341 227 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=6480 $D=0
M1631 348 342 228 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=11110 $D=0
M1632 10 346 966 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=1850 $D=0
M1633 10 347 967 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=6480 $D=0
M1634 10 348 968 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=11110 $D=0
M1635 349 966 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=1850 $D=0
M1636 350 967 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=6480 $D=0
M1637 351 968 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=11110 $D=0
M1638 346 41 349 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=1850 $D=0
M1639 347 41 350 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=6480 $D=0
M1640 348 41 351 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=11110 $D=0
M1641 349 343 241 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=1850 $D=0
M1642 350 344 242 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=6480 $D=0
M1643 351 345 243 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=11110 $D=0
M1644 247 352 349 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=1850 $D=0
M1645 248 353 350 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=6480 $D=0
M1646 249 354 351 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=11110 $D=0
M1647 352 43 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=1850 $D=0
M1648 353 43 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=6480 $D=0
M1649 354 43 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=11110 $D=0
M1650 10 44 355 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=1850 $D=0
M1651 10 44 356 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=6480 $D=0
M1652 10 44 357 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=11110 $D=0
M1653 358 45 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=1850 $D=0
M1654 359 45 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=6480 $D=0
M1655 360 45 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=11110 $D=0
M1656 361 355 226 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=1850 $D=0
M1657 362 356 227 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=6480 $D=0
M1658 363 357 228 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=11110 $D=0
M1659 10 361 969 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=1850 $D=0
M1660 10 362 970 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=6480 $D=0
M1661 10 363 971 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=11110 $D=0
M1662 364 969 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=1850 $D=0
M1663 365 970 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=6480 $D=0
M1664 366 971 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=11110 $D=0
M1665 361 44 364 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=1850 $D=0
M1666 362 44 365 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=6480 $D=0
M1667 363 44 366 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=11110 $D=0
M1668 364 358 241 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=1850 $D=0
M1669 365 359 242 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=6480 $D=0
M1670 366 360 243 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=11110 $D=0
M1671 247 367 364 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=1850 $D=0
M1672 248 368 365 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=6480 $D=0
M1673 249 369 366 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=11110 $D=0
M1674 367 46 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=1850 $D=0
M1675 368 46 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=6480 $D=0
M1676 369 46 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=11110 $D=0
M1677 10 47 370 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=1850 $D=0
M1678 10 47 371 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=6480 $D=0
M1679 10 47 372 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=11110 $D=0
M1680 373 48 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=1850 $D=0
M1681 374 48 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=6480 $D=0
M1682 375 48 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=11110 $D=0
M1683 376 370 226 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=1850 $D=0
M1684 377 371 227 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=6480 $D=0
M1685 378 372 228 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=11110 $D=0
M1686 10 376 972 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=1850 $D=0
M1687 10 377 973 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=6480 $D=0
M1688 10 378 974 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=11110 $D=0
M1689 379 972 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=1850 $D=0
M1690 380 973 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=6480 $D=0
M1691 381 974 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=11110 $D=0
M1692 376 47 379 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=1850 $D=0
M1693 377 47 380 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=6480 $D=0
M1694 378 47 381 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=11110 $D=0
M1695 379 373 241 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=1850 $D=0
M1696 380 374 242 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=6480 $D=0
M1697 381 375 243 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=11110 $D=0
M1698 247 382 379 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=1850 $D=0
M1699 248 383 380 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=6480 $D=0
M1700 249 384 381 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=11110 $D=0
M1701 382 49 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=1850 $D=0
M1702 383 49 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=6480 $D=0
M1703 384 49 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=11110 $D=0
M1704 10 50 385 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=1850 $D=0
M1705 10 50 386 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=6480 $D=0
M1706 10 50 387 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=11110 $D=0
M1707 388 51 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=1850 $D=0
M1708 389 51 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=6480 $D=0
M1709 390 51 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=11110 $D=0
M1710 391 385 226 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=1850 $D=0
M1711 392 386 227 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=6480 $D=0
M1712 393 387 228 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=11110 $D=0
M1713 10 391 975 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=1850 $D=0
M1714 10 392 976 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=6480 $D=0
M1715 10 393 977 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=11110 $D=0
M1716 394 975 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=1850 $D=0
M1717 395 976 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=6480 $D=0
M1718 396 977 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=11110 $D=0
M1719 391 50 394 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=1850 $D=0
M1720 392 50 395 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=6480 $D=0
M1721 393 50 396 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=11110 $D=0
M1722 394 388 241 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=1850 $D=0
M1723 395 389 242 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=6480 $D=0
M1724 396 390 243 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=11110 $D=0
M1725 247 397 394 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=1850 $D=0
M1726 248 398 395 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=6480 $D=0
M1727 249 399 396 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=11110 $D=0
M1728 397 52 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=1850 $D=0
M1729 398 52 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=6480 $D=0
M1730 399 52 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=11110 $D=0
M1731 10 53 400 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=1850 $D=0
M1732 10 53 401 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=6480 $D=0
M1733 10 53 402 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=11110 $D=0
M1734 403 54 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=1850 $D=0
M1735 404 54 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=6480 $D=0
M1736 405 54 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=11110 $D=0
M1737 406 400 226 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=1850 $D=0
M1738 407 401 227 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=6480 $D=0
M1739 408 402 228 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=11110 $D=0
M1740 10 406 978 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=1850 $D=0
M1741 10 407 979 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=6480 $D=0
M1742 10 408 980 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=11110 $D=0
M1743 409 978 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=1850 $D=0
M1744 410 979 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=6480 $D=0
M1745 411 980 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=11110 $D=0
M1746 406 53 409 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=1850 $D=0
M1747 407 53 410 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=6480 $D=0
M1748 408 53 411 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=11110 $D=0
M1749 409 403 241 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=1850 $D=0
M1750 410 404 242 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=6480 $D=0
M1751 411 405 243 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=11110 $D=0
M1752 247 412 409 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=1850 $D=0
M1753 248 413 410 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=6480 $D=0
M1754 249 414 411 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=11110 $D=0
M1755 412 55 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=1850 $D=0
M1756 413 55 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=6480 $D=0
M1757 414 55 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=11110 $D=0
M1758 10 56 415 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=1850 $D=0
M1759 10 56 416 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=6480 $D=0
M1760 10 56 417 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=11110 $D=0
M1761 418 57 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=1850 $D=0
M1762 419 57 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=6480 $D=0
M1763 420 57 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=11110 $D=0
M1764 421 415 226 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=1850 $D=0
M1765 422 416 227 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=6480 $D=0
M1766 423 417 228 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=11110 $D=0
M1767 10 421 981 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=1850 $D=0
M1768 10 422 982 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=6480 $D=0
M1769 10 423 983 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=11110 $D=0
M1770 424 981 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=1850 $D=0
M1771 425 982 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=6480 $D=0
M1772 426 983 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=11110 $D=0
M1773 421 56 424 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=1850 $D=0
M1774 422 56 425 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=6480 $D=0
M1775 423 56 426 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=11110 $D=0
M1776 424 418 241 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=1850 $D=0
M1777 425 419 242 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=6480 $D=0
M1778 426 420 243 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=11110 $D=0
M1779 247 427 424 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=1850 $D=0
M1780 248 428 425 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=6480 $D=0
M1781 249 429 426 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=11110 $D=0
M1782 427 58 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=1850 $D=0
M1783 428 58 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=6480 $D=0
M1784 429 58 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=11110 $D=0
M1785 10 59 430 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=1850 $D=0
M1786 10 59 431 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=6480 $D=0
M1787 10 59 432 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=11110 $D=0
M1788 433 60 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=1850 $D=0
M1789 434 60 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=6480 $D=0
M1790 435 60 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=11110 $D=0
M1791 436 430 226 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=1850 $D=0
M1792 437 431 227 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=6480 $D=0
M1793 438 432 228 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=11110 $D=0
M1794 10 436 984 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=1850 $D=0
M1795 10 437 985 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=6480 $D=0
M1796 10 438 986 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=11110 $D=0
M1797 439 984 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=1850 $D=0
M1798 440 985 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=6480 $D=0
M1799 441 986 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=11110 $D=0
M1800 436 59 439 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=1850 $D=0
M1801 437 59 440 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=6480 $D=0
M1802 438 59 441 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=11110 $D=0
M1803 439 433 241 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=1850 $D=0
M1804 440 434 242 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=6480 $D=0
M1805 441 435 243 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=11110 $D=0
M1806 247 442 439 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=1850 $D=0
M1807 248 443 440 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=6480 $D=0
M1808 249 444 441 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=11110 $D=0
M1809 442 61 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=1850 $D=0
M1810 443 61 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=6480 $D=0
M1811 444 61 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=11110 $D=0
M1812 10 62 445 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=1850 $D=0
M1813 10 62 446 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=6480 $D=0
M1814 10 62 447 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=11110 $D=0
M1815 448 63 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=1850 $D=0
M1816 449 63 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=6480 $D=0
M1817 450 63 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=11110 $D=0
M1818 451 445 226 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=1850 $D=0
M1819 452 446 227 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=6480 $D=0
M1820 453 447 228 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=11110 $D=0
M1821 10 451 987 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=1850 $D=0
M1822 10 452 988 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=6480 $D=0
M1823 10 453 989 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=11110 $D=0
M1824 454 987 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=1850 $D=0
M1825 455 988 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=6480 $D=0
M1826 456 989 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=11110 $D=0
M1827 451 62 454 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=1850 $D=0
M1828 452 62 455 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=6480 $D=0
M1829 453 62 456 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=11110 $D=0
M1830 454 448 241 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=1850 $D=0
M1831 455 449 242 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=6480 $D=0
M1832 456 450 243 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=11110 $D=0
M1833 247 457 454 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=1850 $D=0
M1834 248 458 455 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=6480 $D=0
M1835 249 459 456 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=11110 $D=0
M1836 457 64 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=1850 $D=0
M1837 458 64 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=6480 $D=0
M1838 459 64 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=11110 $D=0
M1839 10 65 460 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=1850 $D=0
M1840 10 65 461 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=6480 $D=0
M1841 10 65 462 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=11110 $D=0
M1842 463 66 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=1850 $D=0
M1843 464 66 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=6480 $D=0
M1844 465 66 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=11110 $D=0
M1845 466 460 226 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=1850 $D=0
M1846 467 461 227 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=6480 $D=0
M1847 468 462 228 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=11110 $D=0
M1848 10 466 990 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=1850 $D=0
M1849 10 467 991 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=6480 $D=0
M1850 10 468 992 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=11110 $D=0
M1851 469 990 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=1850 $D=0
M1852 470 991 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=6480 $D=0
M1853 471 992 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=11110 $D=0
M1854 466 65 469 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=1850 $D=0
M1855 467 65 470 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=6480 $D=0
M1856 468 65 471 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=11110 $D=0
M1857 469 463 241 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=1850 $D=0
M1858 470 464 242 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=6480 $D=0
M1859 471 465 243 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=11110 $D=0
M1860 247 472 469 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=1850 $D=0
M1861 248 473 470 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=6480 $D=0
M1862 249 474 471 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=11110 $D=0
M1863 472 67 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=1850 $D=0
M1864 473 67 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=6480 $D=0
M1865 474 67 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=11110 $D=0
M1866 10 68 475 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=1850 $D=0
M1867 10 68 476 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=6480 $D=0
M1868 10 68 477 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=11110 $D=0
M1869 478 69 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=1850 $D=0
M1870 479 69 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=6480 $D=0
M1871 480 69 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=11110 $D=0
M1872 481 475 226 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=1850 $D=0
M1873 482 476 227 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=6480 $D=0
M1874 483 477 228 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=11110 $D=0
M1875 10 481 993 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=1850 $D=0
M1876 10 482 994 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=6480 $D=0
M1877 10 483 995 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=11110 $D=0
M1878 484 993 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=1850 $D=0
M1879 485 994 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=6480 $D=0
M1880 486 995 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=11110 $D=0
M1881 481 68 484 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=1850 $D=0
M1882 482 68 485 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=6480 $D=0
M1883 483 68 486 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=11110 $D=0
M1884 484 478 241 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=1850 $D=0
M1885 485 479 242 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=6480 $D=0
M1886 486 480 243 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=11110 $D=0
M1887 247 487 484 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=1850 $D=0
M1888 248 488 485 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=6480 $D=0
M1889 249 489 486 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=11110 $D=0
M1890 487 70 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=1850 $D=0
M1891 488 70 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=6480 $D=0
M1892 489 70 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=11110 $D=0
M1893 10 71 490 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=1850 $D=0
M1894 10 71 491 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=6480 $D=0
M1895 10 71 492 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=11110 $D=0
M1896 493 72 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=1850 $D=0
M1897 494 72 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=6480 $D=0
M1898 495 72 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=11110 $D=0
M1899 496 490 226 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=1850 $D=0
M1900 497 491 227 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=6480 $D=0
M1901 498 492 228 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=11110 $D=0
M1902 10 496 996 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=1850 $D=0
M1903 10 497 997 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=6480 $D=0
M1904 10 498 998 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=11110 $D=0
M1905 499 996 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=1850 $D=0
M1906 500 997 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=6480 $D=0
M1907 501 998 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=11110 $D=0
M1908 496 71 499 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=1850 $D=0
M1909 497 71 500 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=6480 $D=0
M1910 498 71 501 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=11110 $D=0
M1911 499 493 241 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=1850 $D=0
M1912 500 494 242 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=6480 $D=0
M1913 501 495 243 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=11110 $D=0
M1914 247 502 499 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=1850 $D=0
M1915 248 503 500 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=6480 $D=0
M1916 249 504 501 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=11110 $D=0
M1917 502 73 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=1850 $D=0
M1918 503 73 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=6480 $D=0
M1919 504 73 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=11110 $D=0
M1920 10 74 505 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=1850 $D=0
M1921 10 74 506 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=6480 $D=0
M1922 10 74 507 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=11110 $D=0
M1923 508 75 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=1850 $D=0
M1924 509 75 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=6480 $D=0
M1925 510 75 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=11110 $D=0
M1926 511 505 226 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=1850 $D=0
M1927 512 506 227 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=6480 $D=0
M1928 513 507 228 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=11110 $D=0
M1929 10 511 999 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=1850 $D=0
M1930 10 512 1000 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=6480 $D=0
M1931 10 513 1001 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=11110 $D=0
M1932 514 999 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=1850 $D=0
M1933 515 1000 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=6480 $D=0
M1934 516 1001 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=11110 $D=0
M1935 511 74 514 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=1850 $D=0
M1936 512 74 515 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=6480 $D=0
M1937 513 74 516 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=11110 $D=0
M1938 514 508 241 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=1850 $D=0
M1939 515 509 242 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=6480 $D=0
M1940 516 510 243 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=11110 $D=0
M1941 247 517 514 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=1850 $D=0
M1942 248 518 515 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=6480 $D=0
M1943 249 519 516 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=11110 $D=0
M1944 517 76 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=1850 $D=0
M1945 518 76 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=6480 $D=0
M1946 519 76 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=11110 $D=0
M1947 10 77 520 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=1850 $D=0
M1948 10 77 521 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=6480 $D=0
M1949 10 77 522 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=11110 $D=0
M1950 523 78 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=1850 $D=0
M1951 524 78 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=6480 $D=0
M1952 525 78 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=11110 $D=0
M1953 526 520 226 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=1850 $D=0
M1954 527 521 227 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=6480 $D=0
M1955 528 522 228 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=11110 $D=0
M1956 10 526 1002 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=1850 $D=0
M1957 10 527 1003 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=6480 $D=0
M1958 10 528 1004 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=11110 $D=0
M1959 529 1002 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=1850 $D=0
M1960 530 1003 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=6480 $D=0
M1961 531 1004 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=11110 $D=0
M1962 526 77 529 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=1850 $D=0
M1963 527 77 530 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=6480 $D=0
M1964 528 77 531 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=11110 $D=0
M1965 529 523 241 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=1850 $D=0
M1966 530 524 242 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=6480 $D=0
M1967 531 525 243 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=11110 $D=0
M1968 247 532 529 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=1850 $D=0
M1969 248 533 530 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=6480 $D=0
M1970 249 534 531 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=11110 $D=0
M1971 532 79 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=1850 $D=0
M1972 533 79 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=6480 $D=0
M1973 534 79 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=11110 $D=0
M1974 10 80 535 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=1850 $D=0
M1975 10 80 536 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=6480 $D=0
M1976 10 80 537 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=11110 $D=0
M1977 538 81 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=1850 $D=0
M1978 539 81 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=6480 $D=0
M1979 540 81 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=11110 $D=0
M1980 541 535 226 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=1850 $D=0
M1981 542 536 227 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=6480 $D=0
M1982 543 537 228 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=11110 $D=0
M1983 10 541 1005 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=1850 $D=0
M1984 10 542 1006 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=6480 $D=0
M1985 10 543 1007 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=11110 $D=0
M1986 544 1005 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=1850 $D=0
M1987 545 1006 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=6480 $D=0
M1988 546 1007 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=11110 $D=0
M1989 541 80 544 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=1850 $D=0
M1990 542 80 545 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=6480 $D=0
M1991 543 80 546 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=11110 $D=0
M1992 544 538 241 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=1850 $D=0
M1993 545 539 242 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=6480 $D=0
M1994 546 540 243 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=11110 $D=0
M1995 247 547 544 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=1850 $D=0
M1996 248 548 545 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=6480 $D=0
M1997 249 549 546 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=11110 $D=0
M1998 547 82 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=1850 $D=0
M1999 548 82 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=6480 $D=0
M2000 549 82 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=11110 $D=0
M2001 10 83 550 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=1850 $D=0
M2002 10 83 551 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=6480 $D=0
M2003 10 83 552 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=11110 $D=0
M2004 553 84 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=1850 $D=0
M2005 554 84 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=6480 $D=0
M2006 555 84 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=11110 $D=0
M2007 556 550 226 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=1850 $D=0
M2008 557 551 227 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=6480 $D=0
M2009 558 552 228 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=11110 $D=0
M2010 10 556 1008 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=1850 $D=0
M2011 10 557 1009 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=6480 $D=0
M2012 10 558 1010 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=11110 $D=0
M2013 559 1008 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=1850 $D=0
M2014 560 1009 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=6480 $D=0
M2015 561 1010 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=11110 $D=0
M2016 556 83 559 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=1850 $D=0
M2017 557 83 560 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=6480 $D=0
M2018 558 83 561 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=11110 $D=0
M2019 559 553 241 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=1850 $D=0
M2020 560 554 242 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=6480 $D=0
M2021 561 555 243 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=11110 $D=0
M2022 247 562 559 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=1850 $D=0
M2023 248 563 560 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=6480 $D=0
M2024 249 564 561 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=11110 $D=0
M2025 562 85 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=1850 $D=0
M2026 563 85 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=6480 $D=0
M2027 564 85 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=11110 $D=0
M2028 10 86 565 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=1850 $D=0
M2029 10 86 566 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=6480 $D=0
M2030 10 86 567 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=11110 $D=0
M2031 568 87 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=1850 $D=0
M2032 569 87 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=6480 $D=0
M2033 570 87 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=11110 $D=0
M2034 571 565 226 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=1850 $D=0
M2035 572 566 227 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=6480 $D=0
M2036 573 567 228 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=11110 $D=0
M2037 10 571 1011 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=1850 $D=0
M2038 10 572 1012 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=6480 $D=0
M2039 10 573 1013 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=11110 $D=0
M2040 574 1011 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=1850 $D=0
M2041 575 1012 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=6480 $D=0
M2042 576 1013 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=11110 $D=0
M2043 571 86 574 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=1850 $D=0
M2044 572 86 575 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=6480 $D=0
M2045 573 86 576 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=11110 $D=0
M2046 574 568 241 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=1850 $D=0
M2047 575 569 242 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=6480 $D=0
M2048 576 570 243 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=11110 $D=0
M2049 247 577 574 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=1850 $D=0
M2050 248 578 575 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=6480 $D=0
M2051 249 579 576 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=11110 $D=0
M2052 577 88 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=1850 $D=0
M2053 578 88 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=6480 $D=0
M2054 579 88 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=11110 $D=0
M2055 10 89 580 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=1850 $D=0
M2056 10 89 581 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=6480 $D=0
M2057 10 89 582 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=11110 $D=0
M2058 583 90 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=1850 $D=0
M2059 584 90 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=6480 $D=0
M2060 585 90 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=11110 $D=0
M2061 586 580 226 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=1850 $D=0
M2062 587 581 227 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=6480 $D=0
M2063 588 582 228 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=11110 $D=0
M2064 10 586 1014 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=1850 $D=0
M2065 10 587 1015 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=6480 $D=0
M2066 10 588 1016 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=11110 $D=0
M2067 589 1014 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=1850 $D=0
M2068 590 1015 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=6480 $D=0
M2069 591 1016 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=11110 $D=0
M2070 586 89 589 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=1850 $D=0
M2071 587 89 590 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=6480 $D=0
M2072 588 89 591 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=11110 $D=0
M2073 589 583 241 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=1850 $D=0
M2074 590 584 242 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=6480 $D=0
M2075 591 585 243 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=11110 $D=0
M2076 247 592 589 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=1850 $D=0
M2077 248 593 590 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=6480 $D=0
M2078 249 594 591 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=11110 $D=0
M2079 592 91 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=1850 $D=0
M2080 593 91 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=6480 $D=0
M2081 594 91 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=11110 $D=0
M2082 10 92 595 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=1850 $D=0
M2083 10 92 596 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=6480 $D=0
M2084 10 92 597 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=11110 $D=0
M2085 598 93 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=1850 $D=0
M2086 599 93 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=6480 $D=0
M2087 600 93 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=11110 $D=0
M2088 601 595 226 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=1850 $D=0
M2089 602 596 227 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=6480 $D=0
M2090 603 597 228 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=11110 $D=0
M2091 10 601 1017 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=1850 $D=0
M2092 10 602 1018 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=6480 $D=0
M2093 10 603 1019 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=11110 $D=0
M2094 604 1017 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=1850 $D=0
M2095 605 1018 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=6480 $D=0
M2096 606 1019 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=11110 $D=0
M2097 601 92 604 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=1850 $D=0
M2098 602 92 605 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=6480 $D=0
M2099 603 92 606 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=11110 $D=0
M2100 604 598 241 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=1850 $D=0
M2101 605 599 242 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=6480 $D=0
M2102 606 600 243 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=11110 $D=0
M2103 247 607 604 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=1850 $D=0
M2104 248 608 605 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=6480 $D=0
M2105 249 609 606 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=11110 $D=0
M2106 607 94 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=1850 $D=0
M2107 608 94 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=6480 $D=0
M2108 609 94 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=11110 $D=0
M2109 10 95 610 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=1850 $D=0
M2110 10 95 611 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=6480 $D=0
M2111 10 95 612 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=11110 $D=0
M2112 613 96 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=1850 $D=0
M2113 614 96 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=6480 $D=0
M2114 615 96 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=11110 $D=0
M2115 616 610 226 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=1850 $D=0
M2116 617 611 227 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=6480 $D=0
M2117 618 612 228 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=11110 $D=0
M2118 10 616 1020 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=1850 $D=0
M2119 10 617 1021 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=6480 $D=0
M2120 10 618 1022 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=11110 $D=0
M2121 619 1020 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=1850 $D=0
M2122 620 1021 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=6480 $D=0
M2123 621 1022 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=11110 $D=0
M2124 616 95 619 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=1850 $D=0
M2125 617 95 620 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=6480 $D=0
M2126 618 95 621 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=11110 $D=0
M2127 619 613 241 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=1850 $D=0
M2128 620 614 242 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=6480 $D=0
M2129 621 615 243 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=11110 $D=0
M2130 247 622 619 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=1850 $D=0
M2131 248 623 620 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=6480 $D=0
M2132 249 624 621 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=11110 $D=0
M2133 622 97 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=1850 $D=0
M2134 623 97 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=6480 $D=0
M2135 624 97 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=11110 $D=0
M2136 10 98 625 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=1850 $D=0
M2137 10 98 626 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=6480 $D=0
M2138 10 98 627 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=11110 $D=0
M2139 628 99 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=1850 $D=0
M2140 629 99 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=6480 $D=0
M2141 630 99 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=11110 $D=0
M2142 631 625 226 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=1850 $D=0
M2143 632 626 227 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=6480 $D=0
M2144 633 627 228 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=11110 $D=0
M2145 10 631 1023 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=1850 $D=0
M2146 10 632 1024 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=6480 $D=0
M2147 10 633 1025 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=11110 $D=0
M2148 634 1023 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=1850 $D=0
M2149 635 1024 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=6480 $D=0
M2150 636 1025 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=11110 $D=0
M2151 631 98 634 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=1850 $D=0
M2152 632 98 635 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=6480 $D=0
M2153 633 98 636 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=11110 $D=0
M2154 634 628 241 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=1850 $D=0
M2155 635 629 242 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=6480 $D=0
M2156 636 630 243 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=11110 $D=0
M2157 247 637 634 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=1850 $D=0
M2158 248 638 635 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=6480 $D=0
M2159 249 639 636 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=11110 $D=0
M2160 637 100 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=1850 $D=0
M2161 638 100 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=6480 $D=0
M2162 639 100 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=11110 $D=0
M2163 10 101 640 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=1850 $D=0
M2164 10 101 641 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=6480 $D=0
M2165 10 101 642 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=11110 $D=0
M2166 643 102 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=1850 $D=0
M2167 644 102 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=6480 $D=0
M2168 645 102 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=11110 $D=0
M2169 646 640 226 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=1850 $D=0
M2170 647 641 227 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=6480 $D=0
M2171 648 642 228 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=11110 $D=0
M2172 10 646 1026 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=1850 $D=0
M2173 10 647 1027 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=6480 $D=0
M2174 10 648 1028 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=11110 $D=0
M2175 649 1026 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=1850 $D=0
M2176 650 1027 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=6480 $D=0
M2177 651 1028 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=11110 $D=0
M2178 646 101 649 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=1850 $D=0
M2179 647 101 650 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=6480 $D=0
M2180 648 101 651 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=11110 $D=0
M2181 649 643 241 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=1850 $D=0
M2182 650 644 242 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=6480 $D=0
M2183 651 645 243 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=11110 $D=0
M2184 247 652 649 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=1850 $D=0
M2185 248 653 650 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=6480 $D=0
M2186 249 654 651 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=11110 $D=0
M2187 652 103 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=1850 $D=0
M2188 653 103 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=6480 $D=0
M2189 654 103 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=11110 $D=0
M2190 10 104 655 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=1850 $D=0
M2191 10 104 656 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=6480 $D=0
M2192 10 104 657 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=11110 $D=0
M2193 658 105 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=1850 $D=0
M2194 659 105 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=6480 $D=0
M2195 660 105 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=11110 $D=0
M2196 661 655 226 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=1850 $D=0
M2197 662 656 227 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=6480 $D=0
M2198 663 657 228 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=11110 $D=0
M2199 10 661 1029 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=1850 $D=0
M2200 10 662 1030 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=6480 $D=0
M2201 10 663 1031 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=11110 $D=0
M2202 664 1029 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=1850 $D=0
M2203 665 1030 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=6480 $D=0
M2204 666 1031 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=11110 $D=0
M2205 661 104 664 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=1850 $D=0
M2206 662 104 665 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=6480 $D=0
M2207 663 104 666 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=11110 $D=0
M2208 664 658 241 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=1850 $D=0
M2209 665 659 242 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=6480 $D=0
M2210 666 660 243 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=11110 $D=0
M2211 247 667 664 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=1850 $D=0
M2212 248 668 665 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=6480 $D=0
M2213 249 669 666 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=11110 $D=0
M2214 667 106 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=1850 $D=0
M2215 668 106 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=6480 $D=0
M2216 669 106 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=11110 $D=0
M2217 10 107 670 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=1850 $D=0
M2218 10 107 671 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=6480 $D=0
M2219 10 107 672 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=11110 $D=0
M2220 673 108 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=1850 $D=0
M2221 674 108 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=6480 $D=0
M2222 675 108 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=11110 $D=0
M2223 676 670 226 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=1850 $D=0
M2224 677 671 227 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=6480 $D=0
M2225 678 672 228 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=11110 $D=0
M2226 10 676 1032 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=1850 $D=0
M2227 10 677 1033 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=6480 $D=0
M2228 10 678 1034 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=11110 $D=0
M2229 679 1032 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=1850 $D=0
M2230 680 1033 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=6480 $D=0
M2231 681 1034 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=11110 $D=0
M2232 676 107 679 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=1850 $D=0
M2233 677 107 680 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=6480 $D=0
M2234 678 107 681 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=11110 $D=0
M2235 679 673 241 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=1850 $D=0
M2236 680 674 242 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=6480 $D=0
M2237 681 675 243 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=11110 $D=0
M2238 247 682 679 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=1850 $D=0
M2239 248 683 680 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=6480 $D=0
M2240 249 684 681 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=11110 $D=0
M2241 682 111 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=1850 $D=0
M2242 683 111 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=6480 $D=0
M2243 684 111 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=11110 $D=0
M2244 10 112 685 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=1850 $D=0
M2245 10 112 686 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=6480 $D=0
M2246 10 112 687 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=11110 $D=0
M2247 688 113 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=1850 $D=0
M2248 689 113 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=6480 $D=0
M2249 690 113 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=11110 $D=0
M2250 691 685 226 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=1850 $D=0
M2251 692 686 227 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=6480 $D=0
M2252 693 687 228 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=11110 $D=0
M2253 10 691 1035 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=1850 $D=0
M2254 10 692 1036 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=6480 $D=0
M2255 10 693 1037 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=11110 $D=0
M2256 694 1035 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=1850 $D=0
M2257 695 1036 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=6480 $D=0
M2258 696 1037 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=11110 $D=0
M2259 691 112 694 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=1850 $D=0
M2260 692 112 695 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=6480 $D=0
M2261 693 112 696 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=11110 $D=0
M2262 694 688 241 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=1850 $D=0
M2263 695 689 242 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=6480 $D=0
M2264 696 690 243 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=11110 $D=0
M2265 247 697 694 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=1850 $D=0
M2266 248 698 695 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=6480 $D=0
M2267 249 699 696 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=11110 $D=0
M2268 697 116 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=1850 $D=0
M2269 698 116 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=6480 $D=0
M2270 699 116 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=11110 $D=0
M2271 10 117 700 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=1850 $D=0
M2272 10 117 701 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=6480 $D=0
M2273 10 117 702 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=11110 $D=0
M2274 703 118 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=1850 $D=0
M2275 704 118 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=6480 $D=0
M2276 705 118 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=11110 $D=0
M2277 7 703 241 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=1850 $D=0
M2278 7 704 242 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=6480 $D=0
M2279 7 705 243 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=11110 $D=0
M2280 247 700 7 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=1850 $D=0
M2281 248 701 7 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=6480 $D=0
M2282 249 702 7 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=11110 $D=0
M2283 10 709 706 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=1850 $D=0
M2284 10 710 707 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=6480 $D=0
M2285 10 711 708 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=11110 $D=0
M2286 709 119 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=1850 $D=0
M2287 710 119 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=6480 $D=0
M2288 711 119 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=11110 $D=0
M2289 1038 241 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=1850 $D=0
M2290 1039 242 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=6480 $D=0
M2291 1040 243 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=11110 $D=0
M2292 712 709 1038 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=1850 $D=0
M2293 713 710 1039 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=6480 $D=0
M2294 714 711 1040 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=11110 $D=0
M2295 10 712 120 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=1850 $D=0
M2296 10 713 715 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=6480 $D=0
M2297 10 714 716 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=11110 $D=0
M2298 1041 120 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=1850 $D=0
M2299 1042 715 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=6480 $D=0
M2300 1043 716 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=11110 $D=0
M2301 712 706 1041 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=1850 $D=0
M2302 713 707 1042 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=6480 $D=0
M2303 714 708 1043 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=11110 $D=0
M2304 10 720 717 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=1850 $D=0
M2305 10 721 718 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=6480 $D=0
M2306 10 722 719 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=11110 $D=0
M2307 720 119 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=1850 $D=0
M2308 721 119 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=6480 $D=0
M2309 722 119 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=11110 $D=0
M2310 1044 247 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=1850 $D=0
M2311 1045 248 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=6480 $D=0
M2312 1046 249 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=11110 $D=0
M2313 723 720 1044 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=1850 $D=0
M2314 724 721 1045 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=6480 $D=0
M2315 725 722 1046 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=11110 $D=0
M2316 10 723 121 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=1850 $D=0
M2317 10 724 122 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=6480 $D=0
M2318 10 725 123 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=11110 $D=0
M2319 1047 121 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=1850 $D=0
M2320 1048 122 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=6480 $D=0
M2321 1049 123 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=11110 $D=0
M2322 723 717 1047 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=1850 $D=0
M2323 724 718 1048 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=6480 $D=0
M2324 725 719 1049 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=11110 $D=0
M2325 726 124 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=1850 $D=0
M2326 727 124 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=6480 $D=0
M2327 728 124 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=11110 $D=0
M2328 729 124 120 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=1850 $D=0
M2329 730 124 715 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=6480 $D=0
M2330 731 124 716 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=11110 $D=0
M2331 125 726 729 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=1850 $D=0
M2332 126 727 730 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=6480 $D=0
M2333 127 728 731 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=11110 $D=0
M2334 732 128 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=1850 $D=0
M2335 733 128 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=6480 $D=0
M2336 734 128 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=11110 $D=0
M2337 735 128 121 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=1850 $D=0
M2338 736 128 122 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=6480 $D=0
M2339 737 128 123 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=11110 $D=0
M2340 1050 732 735 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=1850 $D=0
M2341 1051 733 736 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=6480 $D=0
M2342 1052 734 737 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=11110 $D=0
M2343 10 121 1050 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=1850 $D=0
M2344 10 122 1051 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=6480 $D=0
M2345 10 123 1052 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=11110 $D=0
M2346 738 129 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=1850 $D=0
M2347 739 129 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=6480 $D=0
M2348 740 129 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=11110 $D=0
M2349 741 129 735 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=1850 $D=0
M2350 742 129 736 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=6480 $D=0
M2351 743 129 737 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=11110 $D=0
M2352 12 738 741 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=1850 $D=0
M2353 13 739 742 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=6480 $D=0
M2354 14 740 743 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=11110 $D=0
M2355 746 744 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=1850 $D=0
M2356 747 745 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=6480 $D=0
M2357 748 130 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=11110 $D=0
M2358 10 752 749 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=1850 $D=0
M2359 10 753 750 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=6480 $D=0
M2360 10 754 751 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=11110 $D=0
M2361 755 729 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=1850 $D=0
M2362 756 730 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=6480 $D=0
M2363 757 731 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=11110 $D=0
M2364 752 729 744 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=1850 $D=0
M2365 753 730 745 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=6480 $D=0
M2366 754 731 130 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=11110 $D=0
M2367 746 755 752 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=1850 $D=0
M2368 747 756 753 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=6480 $D=0
M2369 748 757 754 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=11110 $D=0
M2370 758 749 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=1850 $D=0
M2371 759 750 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=6480 $D=0
M2372 760 751 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=11110 $D=0
M2373 761 749 741 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=1850 $D=0
M2374 744 750 742 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=6480 $D=0
M2375 745 751 743 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=11110 $D=0
M2376 729 758 761 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=1850 $D=0
M2377 730 759 744 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=6480 $D=0
M2378 731 760 745 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=11110 $D=0
M2379 762 761 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=1850 $D=0
M2380 763 744 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=6480 $D=0
M2381 764 745 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=11110 $D=0
M2382 765 749 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=1850 $D=0
M2383 766 750 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=6480 $D=0
M2384 767 751 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=11110 $D=0
M2385 768 749 762 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=1850 $D=0
M2386 769 750 763 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=6480 $D=0
M2387 770 751 764 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=11110 $D=0
M2388 741 765 768 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=1850 $D=0
M2389 742 766 769 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=6480 $D=0
M2390 743 767 770 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=11110 $D=0
M2391 1068 729 10 10 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=1490 $D=0
M2392 1069 730 10 10 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=6120 $D=0
M2393 1070 731 10 10 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=10750 $D=0
M2394 771 741 1068 10 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=1490 $D=0
M2395 772 742 1069 10 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=6120 $D=0
M2396 773 743 1070 10 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=10750 $D=0
M2397 774 768 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=1850 $D=0
M2398 775 769 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=6480 $D=0
M2399 776 770 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=11110 $D=0
M2400 777 729 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=1850 $D=0
M2401 778 730 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=6480 $D=0
M2402 779 731 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=11110 $D=0
M2403 10 741 777 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=1850 $D=0
M2404 10 742 778 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=6480 $D=0
M2405 10 743 779 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=11110 $D=0
M2406 780 729 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=1850 $D=0
M2407 781 730 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=6480 $D=0
M2408 782 731 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=11110 $D=0
M2409 10 741 780 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=1850 $D=0
M2410 10 742 781 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=6480 $D=0
M2411 10 743 782 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=11110 $D=0
M2412 1071 729 10 10 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=1670 $D=0
M2413 1072 730 10 10 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=6300 $D=0
M2414 1073 731 10 10 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=10930 $D=0
M2415 786 741 1071 10 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=1670 $D=0
M2416 787 742 1072 10 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=6300 $D=0
M2417 788 743 1073 10 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=10930 $D=0
M2418 10 780 786 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=1850 $D=0
M2419 10 781 787 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=6480 $D=0
M2420 10 782 788 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=11110 $D=0
M2421 789 134 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=1850 $D=0
M2422 790 134 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=6480 $D=0
M2423 791 134 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=11110 $D=0
M2424 792 134 771 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=1850 $D=0
M2425 793 134 772 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=6480 $D=0
M2426 794 134 773 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=11110 $D=0
M2427 777 789 792 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=1850 $D=0
M2428 778 790 793 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=6480 $D=0
M2429 779 791 794 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=11110 $D=0
M2430 795 134 774 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=1850 $D=0
M2431 796 134 775 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=6480 $D=0
M2432 797 134 776 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=11110 $D=0
M2433 786 789 795 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=1850 $D=0
M2434 787 790 796 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=6480 $D=0
M2435 788 791 797 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=11110 $D=0
M2436 798 135 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=1850 $D=0
M2437 799 135 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=6480 $D=0
M2438 800 135 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=11110 $D=0
M2439 801 135 795 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=1850 $D=0
M2440 802 135 796 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=6480 $D=0
M2441 803 135 797 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=11110 $D=0
M2442 792 798 801 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=1850 $D=0
M2443 793 799 802 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=6480 $D=0
M2444 794 800 803 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=11110 $D=0
M2445 15 801 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=1850 $D=0
M2446 16 802 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=6480 $D=0
M2447 17 803 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=11110 $D=0
M2448 804 136 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=1850 $D=0
M2449 805 136 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=6480 $D=0
M2450 806 136 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=11110 $D=0
M2451 808 136 807 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=1850 $D=0
M2452 809 136 137 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=6480 $D=0
M2453 810 136 138 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=11110 $D=0
M2454 139 804 808 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=1850 $D=0
M2455 811 805 809 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=6480 $D=0
M2456 807 806 810 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=11110 $D=0
M2457 812 136 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=1850 $D=0
M2458 813 136 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=6480 $D=0
M2459 814 136 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=11110 $D=0
M2460 815 136 140 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=1850 $D=0
M2461 816 136 141 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=6480 $D=0
M2462 817 136 142 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=11110 $D=0
M2463 139 812 815 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=1850 $D=0
M2464 139 813 816 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=6480 $D=0
M2465 818 814 817 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=11110 $D=0
M2466 819 136 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=1850 $D=0
M2467 820 136 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=6480 $D=0
M2468 821 136 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=11110 $D=0
M2469 822 136 133 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=1850 $D=0
M2470 823 136 132 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=6480 $D=0
M2471 824 136 131 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=11110 $D=0
M2472 139 819 822 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=1850 $D=0
M2473 139 820 823 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=6480 $D=0
M2474 139 821 824 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=11110 $D=0
M2475 825 136 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=1850 $D=0
M2476 826 136 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=6480 $D=0
M2477 827 136 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=11110 $D=0
M2478 828 136 143 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=1850 $D=0
M2479 829 136 144 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=6480 $D=0
M2480 830 136 145 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=11110 $D=0
M2481 139 825 828 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=1850 $D=0
M2482 139 826 829 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=6480 $D=0
M2483 139 827 830 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=11110 $D=0
M2484 831 136 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=1850 $D=0
M2485 832 136 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=6480 $D=0
M2486 833 136 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=11110 $D=0
M2487 834 136 146 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=1850 $D=0
M2488 835 136 147 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=6480 $D=0
M2489 836 136 148 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=11110 $D=0
M2490 139 831 834 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=1850 $D=0
M2491 139 832 835 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=6480 $D=0
M2492 139 833 836 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=11110 $D=0
M2493 10 729 1053 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=1850 $D=0
M2494 10 730 1054 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=6480 $D=0
M2495 10 731 1055 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=11110 $D=0
M2496 811 1053 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=1850 $D=0
M2497 807 1054 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=6480 $D=0
M2498 137 1055 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=11110 $D=0
M2499 837 149 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=1850 $D=0
M2500 838 149 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=6480 $D=0
M2501 839 149 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=11110 $D=0
M2502 818 149 811 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=1850 $D=0
M2503 150 149 807 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=6480 $D=0
M2504 140 149 137 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=11110 $D=0
M2505 808 837 818 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=1850 $D=0
M2506 809 838 150 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=6480 $D=0
M2507 810 839 140 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=11110 $D=0
M2508 840 151 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=1850 $D=0
M2509 841 151 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=6480 $D=0
M2510 842 151 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=11110 $D=0
M2511 152 151 818 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=1850 $D=0
M2512 153 151 150 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=6480 $D=0
M2513 154 151 140 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=11110 $D=0
M2514 815 840 152 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=1850 $D=0
M2515 816 841 153 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=6480 $D=0
M2516 817 842 154 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=11110 $D=0
M2517 843 155 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=1850 $D=0
M2518 844 155 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=6480 $D=0
M2519 845 155 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=11110 $D=0
M2520 110 155 152 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=1850 $D=0
M2521 114 155 153 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=6480 $D=0
M2522 109 155 154 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=11110 $D=0
M2523 822 843 110 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=1850 $D=0
M2524 823 844 114 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=6480 $D=0
M2525 824 845 109 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=11110 $D=0
M2526 846 156 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=1850 $D=0
M2527 847 156 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=6480 $D=0
M2528 848 156 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=11110 $D=0
M2529 157 156 110 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=1850 $D=0
M2530 158 156 114 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=6480 $D=0
M2531 159 156 109 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=11110 $D=0
M2532 828 846 157 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=1850 $D=0
M2533 829 847 158 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=6480 $D=0
M2534 830 848 159 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=11110 $D=0
M2535 849 160 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=1850 $D=0
M2536 850 160 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=6480 $D=0
M2537 851 160 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=11110 $D=0
M2538 205 160 157 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=1850 $D=0
M2539 206 160 158 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=6480 $D=0
M2540 207 160 159 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=11110 $D=0
M2541 834 849 205 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=1850 $D=0
M2542 835 850 206 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=6480 $D=0
M2543 836 851 207 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=11110 $D=0
M2544 852 161 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=1850 $D=0
M2545 853 161 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=6480 $D=0
M2546 854 161 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=11110 $D=0
M2547 162 161 121 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=1850 $D=0
M2548 855 161 122 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=6480 $D=0
M2549 856 161 123 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=11110 $D=0
M2550 12 852 162 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=1850 $D=0
M2551 13 853 855 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=6480 $D=0
M2552 14 854 856 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=11110 $D=0
M2553 857 120 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=1850 $D=0
M2554 858 715 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=6480 $D=0
M2555 859 716 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=11110 $D=0
M2556 10 162 857 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=1850 $D=0
M2557 10 855 858 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=6480 $D=0
M2558 10 856 859 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=11110 $D=0
M2559 1074 120 10 10 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=1670 $D=0
M2560 1075 715 10 10 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=6300 $D=0
M2561 1076 716 10 10 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=10930 $D=0
M2562 863 162 1074 10 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=1670 $D=0
M2563 864 855 1075 10 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=6300 $D=0
M2564 865 856 1076 10 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=10930 $D=0
M2565 10 857 863 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=1850 $D=0
M2566 10 858 864 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=6480 $D=0
M2567 10 859 865 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=11110 $D=0
M2568 1056 10 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=1850 $D=0
M2569 1057 866 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=6480 $D=0
M2570 1058 867 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=11110 $D=0
M2571 10 863 1056 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=1850 $D=0
M2572 10 864 1057 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=6480 $D=0
M2573 10 865 1058 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=11110 $D=0
M2574 866 1056 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=1850 $D=0
M2575 867 1057 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=6480 $D=0
M2576 163 1058 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=11110 $D=0
M2577 1077 120 10 10 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=1490 $D=0
M2578 1078 715 10 10 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=6120 $D=0
M2579 1079 716 10 10 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=10750 $D=0
M2580 868 871 1077 10 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=1490 $D=0
M2581 869 872 1078 10 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=6120 $D=0
M2582 870 873 1079 10 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=10750 $D=0
M2583 871 162 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=1850 $D=0
M2584 872 855 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=6480 $D=0
M2585 873 856 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=11110 $D=0
M2586 874 868 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=1850 $D=0
M2587 875 869 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=6480 $D=0
M2588 876 870 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=11110 $D=0
M2589 10 10 874 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=1850 $D=0
M2590 10 866 875 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=6480 $D=0
M2591 10 867 876 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=11110 $D=0
M2592 879 7 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=1850 $D=0
M2593 880 877 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=6480 $D=0
M2594 881 878 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=11110 $D=0
M2595 877 874 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=1850 $D=0
M2596 878 875 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=6480 $D=0
M2597 164 876 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=11110 $D=0
M2598 10 879 877 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=1850 $D=0
M2599 10 880 878 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=6480 $D=0
M2600 10 881 164 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=11110 $D=0
M2601 884 882 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=1850 $D=0
M2602 885 883 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=6480 $D=0
M2603 886 165 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=11110 $D=0
M2604 10 890 887 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=1850 $D=0
M2605 10 891 888 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=6480 $D=0
M2606 10 892 889 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=11110 $D=0
M2607 893 125 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=1850 $D=0
M2608 894 126 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=6480 $D=0
M2609 895 127 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=11110 $D=0
M2610 890 125 882 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=1850 $D=0
M2611 891 126 883 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=6480 $D=0
M2612 892 127 165 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=11110 $D=0
M2613 884 893 890 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=1850 $D=0
M2614 885 894 891 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=6480 $D=0
M2615 886 895 892 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=11110 $D=0
M2616 896 887 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=1850 $D=0
M2617 897 888 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=6480 $D=0
M2618 898 889 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=11110 $D=0
M2619 899 887 7 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=1850 $D=0
M2620 882 888 7 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=6480 $D=0
M2621 883 889 7 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=11110 $D=0
M2622 125 896 899 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=1850 $D=0
M2623 126 897 882 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=6480 $D=0
M2624 127 898 883 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=11110 $D=0
M2625 900 899 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=1850 $D=0
M2626 901 882 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=6480 $D=0
M2627 902 883 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=11110 $D=0
M2628 903 887 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=1850 $D=0
M2629 904 888 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=6480 $D=0
M2630 905 889 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=11110 $D=0
M2631 208 887 900 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=1850 $D=0
M2632 209 888 901 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=6480 $D=0
M2633 210 889 902 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=11110 $D=0
M2634 7 903 208 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=1850 $D=0
M2635 7 904 209 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=6480 $D=0
M2636 7 905 210 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=11110 $D=0
M2637 906 166 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=1850 $D=0
M2638 907 166 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=6480 $D=0
M2639 908 166 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=11110 $D=0
M2640 909 166 208 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=1850 $D=0
M2641 910 166 209 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=6480 $D=0
M2642 911 166 210 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=11110 $D=0
M2643 15 906 909 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=1850 $D=0
M2644 16 907 910 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=6480 $D=0
M2645 17 908 911 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=11110 $D=0
M2646 912 167 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=1850 $D=0
M2647 913 167 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=6480 $D=0
M2648 914 167 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=11110 $D=0
M2649 915 167 909 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=1850 $D=0
M2650 916 167 910 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=6480 $D=0
M2651 917 167 911 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=11110 $D=0
M2652 7 912 915 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=1850 $D=0
M2653 10 913 916 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=6480 $D=0
M2654 10 914 917 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=11110 $D=0
M2655 918 119 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=1850 $D=0
M2656 919 119 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=6480 $D=0
M2657 920 119 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=11110 $D=0
M2658 10 918 921 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=1850 $D=0
M2659 10 919 922 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=6480 $D=0
M2660 10 920 923 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=11110 $D=0
M2661 924 119 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=1850 $D=0
M2662 925 119 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=6480 $D=0
M2663 926 119 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=11110 $D=0
M2664 927 921 915 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=1850 $D=0
M2665 928 922 916 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=6480 $D=0
M2666 929 923 917 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=11110 $D=0
M2667 10 927 1059 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=1850 $D=0
M2668 10 928 1060 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=6480 $D=0
M2669 10 929 1061 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=11110 $D=0
M2670 930 1059 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=1850 $D=0
M2671 931 1060 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=6480 $D=0
M2672 932 1061 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=11110 $D=0
M2673 927 918 930 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=1850 $D=0
M2674 928 919 931 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=6480 $D=0
M2675 929 920 932 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=11110 $D=0
M2676 933 924 930 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=1850 $D=0
M2677 934 925 931 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=6480 $D=0
M2678 935 926 932 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=11110 $D=0
M2679 10 939 936 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=1850 $D=0
M2680 10 940 937 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=6480 $D=0
M2681 10 941 938 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=11110 $D=0
M2682 939 119 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=1850 $D=0
M2683 940 119 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=6480 $D=0
M2684 941 119 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=11110 $D=0
M2685 1062 933 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=1850 $D=0
M2686 1063 934 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=6480 $D=0
M2687 1064 935 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=11110 $D=0
M2688 942 939 1062 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=1850 $D=0
M2689 943 940 1063 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=6480 $D=0
M2690 944 941 1064 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=11110 $D=0
M2691 10 942 125 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=1850 $D=0
M2692 10 943 126 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=6480 $D=0
M2693 10 944 127 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=11110 $D=0
M2694 1065 125 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=1850 $D=0
M2695 1066 126 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=6480 $D=0
M2696 1067 127 10 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=11110 $D=0
M2697 942 936 1065 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=1850 $D=0
M2698 943 937 1066 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=6480 $D=0
M2699 944 938 1067 10 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=11110 $D=0
.ENDS
***************************************
.SUBCKT datapath vss! vdd! mem_mux_sel<0> dmem_rdata<2> dmem_rdata<1> dmem_rdata<0> mem_mux_sel<1> mem_mux_sel<2> rd_mux_sel<0> cmp_out imm<2> imm<1> imm<0> rd_mux_sel<1> rd_mux_sel<2> rd_sel<31> rs1_sel<31> rs2_sel<31> rd_sel<30> rs1_sel<30>
+ rs2_sel<30> rd_sel<29> rs1_sel<29> rs2_sel<29> rd_sel<28> rs1_sel<28> rs2_sel<28> rd_sel<27> rs1_sel<27> rs2_sel<27> rd_sel<26> rs1_sel<26> rs2_sel<26> rd_sel<25> rs1_sel<25> rs2_sel<25> rd_sel<24> rs1_sel<24> rs2_sel<24> rd_sel<23>
+ rs1_sel<23> rs2_sel<23> rd_sel<22> rs1_sel<22> rs2_sel<22> rd_sel<21> rs1_sel<21> rs2_sel<21> rd_sel<20> rs1_sel<20> rs2_sel<20> rd_sel<19> rs1_sel<19> rs2_sel<19> rd_sel<18> rs1_sel<18> rs2_sel<18> rd_sel<17> rs1_sel<17> rs2_sel<17>
+ rd_sel<16> rs1_sel<16> rs2_sel<16> rd_sel<15> rs1_sel<15> rs2_sel<15> rd_sel<14> rs1_sel<14> rs2_sel<14> rd_sel<13> rs1_sel<13> rs2_sel<13> rd_sel<12> rs1_sel<12> rs2_sel<12> rd_sel<11> rs1_sel<11> rs2_sel<11> rd_sel<10> rs1_sel<10>
+ rs2_sel<10> rd_sel<9> rs1_sel<9> rs2_sel<9> rd_sel<8> rs1_sel<8> rs2_sel<8> rd_sel<7> rs1_sel<7> rs2_sel<7> rd_sel<6> rs1_sel<6> rs2_sel<6> rd_sel<5> rs1_sel<5> rs2_sel<5> rd_sel<4> rs1_sel<4> rs2_sel<4> rd_sel<3>
+ rs1_sel<3> rs2_sel<3> rd_sel<2> rs1_sel<2> rs2_sel<2> rd_sel<1> rs1_sel<1> rs2_sel<1> rs2_sel<0> rs1_sel<0> clk dmem_wdata<2> dmem_wdata<1> dmem_wdata<0> alu_mux_1_sel alu_inv_rs2 alu_mux_2_sel alu_cin alu_op<0> alu_op<1>
+ dmem_addr<2> dmem_addr<1> dmem_addr<0> shift_dir cmp_mux_sel cmp_eq cmp_lt pc_mux_sel rst imem_addr<2> imem_addr<1> imem_addr<0> dmem_rdata<4> dmem_rdata<3> imm<4> imm<3> dmem_wdata<4> dmem_wdata<3> dmem_addr<3> dmem_addr<4>
+ imem_addr<4> imem_addr<3> dmem_rdata<6> dmem_rdata<5> imm<6> imm<5> dmem_wdata<6> dmem_wdata<5> dmem_addr<6> dmem_addr<5> imem_addr<6> imem_addr<5> dmem_rdata<8> dmem_rdata<7> imm<8> imm<7> dmem_wdata<8> dmem_wdata<7> dmem_addr<8> dmem_addr<7>
+ imem_addr<8> imem_addr<7> dmem_rdata<10> dmem_rdata<9> imm<10> imm<9> dmem_wdata<10> dmem_wdata<9> dmem_addr<9> dmem_addr<10> imem_addr<10> imem_addr<9> dmem_rdata<12> dmem_rdata<11> imm<12> imm<11> dmem_wdata<12> dmem_wdata<11> dmem_addr<11> dmem_addr<12>
+ imem_addr<12> imem_addr<11> dmem_rdata<14> dmem_rdata<13> imm<14> imm<13> dmem_wdata<14> dmem_wdata<13> dmem_addr<14> dmem_addr<13> imem_addr<14> imem_addr<13> dmem_rdata<16> dmem_rdata<15> imm<16> imm<15> dmem_wdata<16> dmem_wdata<15> dmem_addr<16> dmem_addr<15>
+ shift_msb imem_addr<16> imem_addr<15> dmem_rdata<20> dmem_rdata<19> dmem_rdata<18> dmem_rdata<17> imm<20> imm<19> imm<18> imm<17> dmem_wdata<20> dmem_wdata<19> dmem_wdata<18> dmem_wdata<17> dmem_addr<17> dmem_addr<20> dmem_addr<19> dmem_addr<18> imem_addr<20>
+ imem_addr<19> imem_addr<18> imem_addr<17> dmem_rdata<22> dmem_rdata<21> imm<22> imm<21> dmem_wdata<22> dmem_wdata<21> dmem_addr<22> dmem_addr<21> imem_addr<22> imem_addr<21> dmem_rdata<24> dmem_rdata<23> imm<24> imm<23> dmem_wdata<24> dmem_wdata<23> dmem_addr<24>
+ dmem_addr<23> imem_addr<24> imem_addr<23> dmem_rdata<26> dmem_rdata<25> imm<26> imm<25> dmem_wdata<26> dmem_wdata<25> dmem_addr<26> dmem_addr<25> imem_addr<26> imem_addr<25> dmem_rdata<28> dmem_rdata<27> imm<28> imm<27> dmem_wdata<28> dmem_wdata<27> dmem_addr<28>
+ dmem_addr<27> imem_addr<28> imem_addr<27> dmem_rdata<31> dmem_rdata<30> dmem_rdata<29> imm<31> imm<30> imm<29> dmem_wdata<31> dmem_wdata<30> dmem_wdata<29> dmem_addr<31> dmem_addr<30> dmem_addr<29> cmp_a_31 cmp_b_31 imem_addr<31> imem_addr<30> imem_addr<29>
** N=489 EP=280 IP=2681 FDC=28800
X0 mem_mux_sel<0> dmem_rdata<2> dmem_rdata<1> dmem_rdata<0> mem_mux_sel<1> mem_mux_sel<2> vdd! rd_mux_sel<0> vss! cmp_out imm<2> imm<1> imm<0> dmem_addr<2> dmem_addr<1> dmem_addr<0> rd_mux_sel<1> rd_mux_sel<2> rd_sel<31> rs1_sel<31>
+ rs2_sel<31> rd_sel<30> rs1_sel<30> rs2_sel<30> rd_sel<29> rs1_sel<29> rs2_sel<29> rd_sel<28> rs1_sel<28> rs2_sel<28> rd_sel<27> rs1_sel<27> rs2_sel<27> rd_sel<26> rs1_sel<26> rs2_sel<26> rd_sel<25> rs1_sel<25> rs2_sel<25> rd_sel<24>
+ rs1_sel<24> rs2_sel<24> rd_sel<23> rs1_sel<23> rs2_sel<23> rd_sel<22> rs1_sel<22> rs2_sel<22> rd_sel<21> rs1_sel<21> rs2_sel<21> rd_sel<20> rs1_sel<20> rs2_sel<20> rd_sel<19> rs1_sel<19> rs2_sel<19> rd_sel<18> rs1_sel<18> rs2_sel<18>
+ rd_sel<17> rs1_sel<17> rs2_sel<17> rd_sel<16> rs1_sel<16> rs2_sel<16> rd_sel<15> rs1_sel<15> rs2_sel<15> rd_sel<14> rs1_sel<14> rs2_sel<14> rd_sel<13> rs1_sel<13> rs2_sel<13> rd_sel<12> rs1_sel<12> rs2_sel<12> rd_sel<11> rs1_sel<11>
+ rs2_sel<11> rd_sel<10> rs1_sel<10> rs2_sel<10> rd_sel<9> rs1_sel<9> rs2_sel<9> rd_sel<8> rs1_sel<8> rs2_sel<8> rd_sel<7> rs1_sel<7> rs2_sel<7> rd_sel<6> rs1_sel<6> rs2_sel<6> rd_sel<5> rs1_sel<5> rs2_sel<5> rd_sel<4>
+ rs1_sel<4> rs2_sel<4> rd_sel<3> rs1_sel<3> rs2_sel<3> rd_sel<2> rs1_sel<2> rs2_sel<2> rd_sel<1> rs1_sel<1> rs2_sel<1> rs2_sel<0> rs1_sel<0> clk dmem_wdata<2> dmem_wdata<1> dmem_wdata<0> alu_mux_1_sel imem_addr<2> imem_addr<1>
+ imem_addr<0> alu_inv_rs2 alu_mux_2_sel 153 149 146 alu_cin 129 131 3 132 133 134 135 alu_op<0> alu_op<1> shift_dir 145 143 150
+ 138 151 156 152 160 163 7 147 154 155 148 144 157 167 8 164 158 cmp_mux_sel 161 cmp_eq
+ 165 cmp_lt 168 pc_mux_sel rst
+ ICV_24 $T=0 0 0 0 $X=0 $Y=132400
X1 mem_mux_sel<0> dmem_rdata<4> dmem_rdata<3> mem_mux_sel<1> mem_mux_sel<2> vdd! rd_mux_sel<0> vss! imm<4> imm<3> dmem_addr<4> dmem_addr<3> rd_mux_sel<1> rd_mux_sel<2> rd_sel<31> rs1_sel<31> rs2_sel<31> rd_sel<30> rs1_sel<30> rs2_sel<30>
+ rd_sel<29> rs1_sel<29> rs2_sel<29> rd_sel<28> rs1_sel<28> rs2_sel<28> rd_sel<27> rs1_sel<27> rs2_sel<27> rd_sel<26> rs1_sel<26> rs2_sel<26> rd_sel<25> rs1_sel<25> rs2_sel<25> rd_sel<24> rs1_sel<24> rs2_sel<24> rd_sel<23> rs1_sel<23>
+ rs2_sel<23> rd_sel<22> rs1_sel<22> rs2_sel<22> rd_sel<21> rs1_sel<21> rs2_sel<21> rd_sel<20> rs1_sel<20> rs2_sel<20> rd_sel<19> rs1_sel<19> rs2_sel<19> rd_sel<18> rs1_sel<18> rs2_sel<18> rd_sel<17> rs1_sel<17> rs2_sel<17> rd_sel<16>
+ rs1_sel<16> rs2_sel<16> rd_sel<15> rs1_sel<15> rs2_sel<15> rd_sel<14> rs1_sel<14> rs2_sel<14> rd_sel<13> rs1_sel<13> rs2_sel<13> rd_sel<12> rs1_sel<12> rs2_sel<12> rd_sel<11> rs1_sel<11> rs2_sel<11> rd_sel<10> rs1_sel<10> rs2_sel<10>
+ rd_sel<9> rs1_sel<9> rs2_sel<9> rd_sel<8> rs1_sel<8> rs2_sel<8> rd_sel<7> rs1_sel<7> rs2_sel<7> rd_sel<6> rs1_sel<6> rs2_sel<6> rd_sel<5> rs1_sel<5> rs2_sel<5> rd_sel<4> rs1_sel<4> rs2_sel<4> rd_sel<3> rs1_sel<3>
+ rs2_sel<3> rd_sel<2> rs1_sel<2> rs2_sel<2> rd_sel<1> rs1_sel<1> rs2_sel<1> rs2_sel<0> rs1_sel<0> clk dmem_wdata<4> dmem_wdata<3> alu_mux_1_sel imem_addr<4> imem_addr<3> alu_inv_rs2 alu_mux_2_sel 158 157 129
+ 180 181 4 133 182 alu_op<0> alu_op<1> 183 shift_dir 145 143 188 187 151 144 189 184 191 193 192
+ 194 190 146 150 138 149 160 153 199 198 cmp_mux_sel 195 161 196 165 168 197 pc_mux_sel rst
+ ICV_25 $T=0 0 0 0 $X=0 $Y=123200
X2 mem_mux_sel<0> dmem_rdata<6> dmem_rdata<5> mem_mux_sel<1> mem_mux_sel<2> vdd! rd_mux_sel<0> vss! imm<6> imm<5> dmem_addr<6> dmem_addr<5> rd_mux_sel<1> rd_mux_sel<2> rd_sel<31> rs1_sel<31> rs2_sel<31> rd_sel<30> rs1_sel<30> rs2_sel<30>
+ rd_sel<29> rs1_sel<29> rs2_sel<29> rd_sel<28> rs1_sel<28> rs2_sel<28> rd_sel<27> rs1_sel<27> rs2_sel<27> rd_sel<26> rs1_sel<26> rs2_sel<26> rd_sel<25> rs1_sel<25> rs2_sel<25> rd_sel<24> rs1_sel<24> rs2_sel<24> rd_sel<23> rs1_sel<23>
+ rs2_sel<23> rd_sel<22> rs1_sel<22> rs2_sel<22> rd_sel<21> rs1_sel<21> rs2_sel<21> rd_sel<20> rs1_sel<20> rs2_sel<20> rd_sel<19> rs1_sel<19> rs2_sel<19> rd_sel<18> rs1_sel<18> rs2_sel<18> rd_sel<17> rs1_sel<17> rs2_sel<17> rd_sel<16>
+ rs1_sel<16> rs2_sel<16> rd_sel<15> rs1_sel<15> rs2_sel<15> rd_sel<14> rs1_sel<14> rs2_sel<14> rd_sel<13> rs1_sel<13> rs2_sel<13> rd_sel<12> rs1_sel<12> rs2_sel<12> rd_sel<11> rs1_sel<11> rs2_sel<11> rd_sel<10> rs1_sel<10> rs2_sel<10>
+ rd_sel<9> rs1_sel<9> rs2_sel<9> rd_sel<8> rs1_sel<8> rs2_sel<8> rd_sel<7> rs1_sel<7> rs2_sel<7> rd_sel<6> rs1_sel<6> rs2_sel<6> rd_sel<5> rs1_sel<5> rs2_sel<5> rd_sel<4> rs1_sel<4> rs2_sel<4> rd_sel<3> rs1_sel<3>
+ rs2_sel<3> rd_sel<2> rs1_sel<2> rs2_sel<2> rd_sel<1> rs1_sel<1> rs2_sel<1> rs2_sel<0> rs1_sel<0> clk dmem_wdata<6> dmem_wdata<5> alu_mux_1_sel imem_addr<6> imem_addr<5> alu_inv_rs2 alu_mux_2_sel 180 209 5
+ 208 135 alu_op<0> alu_op<1> shift_dir 188 187 214 213 150 138 215 210 134 219 216 220 217 9 218
+ 146 189 184 149 156 152 153 157 224 225 158 cmp_mux_sel 221 195 222 196 197 223 pc_mux_sel rst
+ ICV_26 $T=0 0 0 0 $X=0 $Y=114000
X3 mem_mux_sel<0> dmem_rdata<8> dmem_rdata<7> vss! mem_mux_sel<1> mem_mux_sel<2> vdd! rd_mux_sel<0> imm<8> imm<7> dmem_addr<8> dmem_addr<7> rd_mux_sel<1> rd_mux_sel<2> rd_sel<31> rs1_sel<31> rs2_sel<31> rd_sel<30> rs1_sel<30> rs2_sel<30>
+ rd_sel<29> rs1_sel<29> rs2_sel<29> rd_sel<28> rs1_sel<28> rs2_sel<28> rd_sel<27> rs1_sel<27> rs2_sel<27> rd_sel<26> rs1_sel<26> rs2_sel<26> rd_sel<25> rs1_sel<25> rs2_sel<25> rd_sel<24> rs1_sel<24> rs2_sel<24> rd_sel<23> rs1_sel<23>
+ rs2_sel<23> rd_sel<22> rs1_sel<22> rs2_sel<22> rd_sel<21> rs1_sel<21> rs2_sel<21> rd_sel<20> rs1_sel<20> rs2_sel<20> rd_sel<19> rs1_sel<19> rs2_sel<19> rd_sel<18> rs1_sel<18> rs2_sel<18> rd_sel<17> rs1_sel<17> rs2_sel<17> rd_sel<16>
+ rs1_sel<16> rs2_sel<16> rd_sel<15> rs1_sel<15> rs2_sel<15> rd_sel<14> rs1_sel<14> rs2_sel<14> rd_sel<13> rs1_sel<13> rs2_sel<13> rd_sel<12> rs1_sel<12> rs2_sel<12> rd_sel<11> rs1_sel<11> rs2_sel<11> rd_sel<10> rs1_sel<10> rs2_sel<10>
+ rd_sel<9> rs1_sel<9> rs2_sel<9> rd_sel<8> rs1_sel<8> rs2_sel<8> rd_sel<7> rs1_sel<7> rs2_sel<7> rd_sel<6> rs1_sel<6> rs2_sel<6> rd_sel<5> rs1_sel<5> rs2_sel<5> rd_sel<4> rs1_sel<4> rs2_sel<4> rd_sel<3> rs1_sel<3>
+ rs2_sel<3> rd_sel<2> rs1_sel<2> rs2_sel<2> rd_sel<1> rs1_sel<1> rs2_sel<1> rs2_sel<0> rs1_sel<0> clk dmem_wdata<8> dmem_wdata<7> alu_mux_1_sel imem_addr<8> imem_addr<7> alu_inv_rs2 234 alu_mux_2_sel 235 208
+ 147 6 237 236 183 alu_op<0> alu_op<1> shift_dir 214 213 242 241 189 184 243 238 160 182 132 244
+ 247 246 146 215 210 149 191 153 157 250 251 158 cmp_mux_sel 245 221 248 222 223 249 pc_mux_sel
+ rst
+ ICV_27 $T=0 0 0 0 $X=0 $Y=104600
X4 mem_mux_sel<0> dmem_rdata<10> dmem_rdata<9> dmem_rdata<7> vss! mem_mux_sel<1> mem_mux_sel<2> vdd! rd_mux_sel<0> imm<10> imm<9> dmem_addr<10> dmem_addr<9> rd_mux_sel<1> rd_mux_sel<2> rd_sel<31> rs1_sel<31> rs2_sel<31> rd_sel<30> rs1_sel<30>
+ rs2_sel<30> rd_sel<29> rs1_sel<29> rs2_sel<29> rd_sel<28> rs1_sel<28> rs2_sel<28> rd_sel<27> rs1_sel<27> rs2_sel<27> rd_sel<26> rs1_sel<26> rs2_sel<26> rd_sel<25> rs1_sel<25> rs2_sel<25> rd_sel<24> rs1_sel<24> rs2_sel<24> rd_sel<23>
+ rs1_sel<23> rs2_sel<23> rd_sel<22> rs1_sel<22> rs2_sel<22> rd_sel<21> rs1_sel<21> rs2_sel<21> rd_sel<20> rs1_sel<20> rs2_sel<20> rd_sel<19> rs1_sel<19> rs2_sel<19> rd_sel<18> rs1_sel<18> rs2_sel<18> rd_sel<17> rs1_sel<17> rs2_sel<17>
+ rd_sel<16> rs1_sel<16> rs2_sel<16> rd_sel<15> rs1_sel<15> rs2_sel<15> rd_sel<14> rs1_sel<14> rs2_sel<14> rd_sel<13> rs1_sel<13> rs2_sel<13> rd_sel<12> rs1_sel<12> rs2_sel<12> rd_sel<11> rs1_sel<11> rs2_sel<11> rd_sel<10> rs1_sel<10>
+ rs2_sel<10> rd_sel<9> rs1_sel<9> rs2_sel<9> rd_sel<8> rs1_sel<8> rs2_sel<8> rd_sel<7> rs1_sel<7> rs2_sel<7> rd_sel<6> rs1_sel<6> rs2_sel<6> rd_sel<5> rs1_sel<5> rs2_sel<5> rd_sel<4> rs1_sel<4> rs2_sel<4> rd_sel<3>
+ rs1_sel<3> rs2_sel<3> rd_sel<2> rs1_sel<2> rs2_sel<2> rd_sel<1> rs1_sel<1> rs2_sel<1> rs2_sel<0> rs1_sel<0> clk dmem_wdata<10> dmem_wdata<9> 260 alu_mux_1_sel 261 imem_addr<10> imem_addr<9> alu_inv_rs2 262
+ 263 alu_mux_2_sel 236 163 7 264 216 alu_op<0> alu_op<1> shift_dir 242 241 269 268 215 210 270 265 156 152
+ 131 3 273 272 146 243 238 149 219 153 157 277 276 158 cmp_mux_sel 271 245 274 248 249
+ 275 pc_mux_sel rst
+ ICV_28 $T=0 0 0 0 $X=0 $Y=95400
X5 mem_mux_sel<0> dmem_rdata<12> dmem_rdata<11> dmem_rdata<7> vss! mem_mux_sel<1> mem_mux_sel<2> vdd! rd_mux_sel<0> imm<12> imm<11> dmem_addr<12> dmem_addr<11> rd_mux_sel<1> rd_mux_sel<2> rd_sel<31> rs1_sel<31> rs2_sel<31> rd_sel<30> rs1_sel<30>
+ rs2_sel<30> rd_sel<29> rs1_sel<29> rs2_sel<29> rd_sel<28> rs1_sel<28> rs2_sel<28> rd_sel<27> rs1_sel<27> rs2_sel<27> rd_sel<26> rs1_sel<26> rs2_sel<26> rd_sel<25> rs1_sel<25> rs2_sel<25> rd_sel<24> rs1_sel<24> rs2_sel<24> rd_sel<23>
+ rs1_sel<23> rs2_sel<23> rd_sel<22> rs1_sel<22> rs2_sel<22> rd_sel<21> rs1_sel<21> rs2_sel<21> rd_sel<20> rs1_sel<20> rs2_sel<20> rd_sel<19> rs1_sel<19> rs2_sel<19> rd_sel<18> rs1_sel<18> rs2_sel<18> rd_sel<17> rs1_sel<17> rs2_sel<17>
+ rd_sel<16> rs1_sel<16> rs2_sel<16> rd_sel<15> rs1_sel<15> rs2_sel<15> rd_sel<14> rs1_sel<14> rs2_sel<14> rd_sel<13> rs1_sel<13> rs2_sel<13> rd_sel<12> rs1_sel<12> rs2_sel<12> rd_sel<11> rs1_sel<11> rs2_sel<11> rd_sel<10> rs1_sel<10>
+ rs2_sel<10> rd_sel<9> rs1_sel<9> rs2_sel<9> rd_sel<8> rs1_sel<8> rs2_sel<8> rd_sel<7> rs1_sel<7> rs2_sel<7> rd_sel<6> rs1_sel<6> rs2_sel<6> rd_sel<5> rs1_sel<5> rs2_sel<5> rd_sel<4> rs1_sel<4> rs2_sel<4> rd_sel<3>
+ rs1_sel<3> rs2_sel<3> rd_sel<2> rs1_sel<2> rs2_sel<2> rd_sel<1> rs1_sel<1> rs2_sel<1> rs2_sel<0> rs1_sel<0> clk dmem_wdata<12> dmem_wdata<11> 286 287 288 289 alu_mux_1_sel imem_addr<12> imem_addr<11>
+ alu_inv_rs2 234 alu_mux_2_sel 264 193 192 290 alu_op<0> alu_op<1> shift_dir 269 268 295 294 243 238 296 291 183 191
+ 181 4 299 298 146 270 265 149 237 153 157 303 302 158 cmp_mux_sel 297 271 300 274 275
+ 301 pc_mux_sel rst
+ ICV_29 $T=0 0 0 0 $X=0 $Y=86200
X6 mem_mux_sel<0> dmem_rdata<14> dmem_rdata<13> dmem_rdata<7> vss! mem_mux_sel<1> mem_mux_sel<2> vdd! rd_mux_sel<0> imm<14> imm<13> dmem_addr<14> dmem_addr<13> rd_mux_sel<1> rd_mux_sel<2> rd_sel<31> rs1_sel<31> rs2_sel<31> rd_sel<30> rs1_sel<30>
+ rs2_sel<30> rd_sel<29> rs1_sel<29> rs2_sel<29> rd_sel<28> rs1_sel<28> rs2_sel<28> rd_sel<27> rs1_sel<27> rs2_sel<27> rd_sel<26> rs1_sel<26> rs2_sel<26> rd_sel<25> rs1_sel<25> rs2_sel<25> rd_sel<24> rs1_sel<24> rs2_sel<24> rd_sel<23>
+ rs1_sel<23> rs2_sel<23> rd_sel<22> rs1_sel<22> rs2_sel<22> rd_sel<21> rs1_sel<21> rs2_sel<21> rd_sel<20> rs1_sel<20> rs2_sel<20> rd_sel<19> rs1_sel<19> rs2_sel<19> rd_sel<18> rs1_sel<18> rs2_sel<18> rd_sel<17> rs1_sel<17> rs2_sel<17>
+ rd_sel<16> rs1_sel<16> rs2_sel<16> rd_sel<15> rs1_sel<15> rs2_sel<15> rd_sel<14> rs1_sel<14> rs2_sel<14> rd_sel<13> rs1_sel<13> rs2_sel<13> rd_sel<12> rs1_sel<12> rs2_sel<12> rd_sel<11> rs1_sel<11> rs2_sel<11> rd_sel<10> rs1_sel<10>
+ rs2_sel<10> rd_sel<9> rs1_sel<9> rs2_sel<9> rd_sel<8> rs1_sel<8> rs2_sel<8> rd_sel<7> rs1_sel<7> rs2_sel<7> rd_sel<6> rs1_sel<6> rs2_sel<6> rd_sel<5> rs1_sel<5> rs2_sel<5> rd_sel<4> rs1_sel<4> rs2_sel<4> rd_sel<3>
+ rs1_sel<3> rs2_sel<3> rd_sel<2> rs1_sel<2> rs2_sel<2> rd_sel<1> rs1_sel<1> rs2_sel<1> rs2_sel<0> rs1_sel<0> clk 220 310 311 312 313 dmem_wdata<14> dmem_wdata<13> alu_mux_1_sel 261
+ imem_addr<14> imem_addr<13> alu_inv_rs2 263 alu_mux_2_sel 290 217 316 alu_op<0> alu_op<1> shift_dir 295 294 321 320 270 265 322 317 219
+ 216 209 5 325 324 146 296 291 149 153 157 329 328 158 cmp_mux_sel 323 297 326 300 301
+ 327 pc_mux_sel rst
+ ICV_30 $T=0 0 0 0 $X=0 $Y=77000
X7 mem_mux_sel<0> dmem_rdata<16> dmem_rdata<15> dmem_rdata<7> vss! mem_mux_sel<1> mem_mux_sel<2> vdd! rd_mux_sel<0> imm<16> imm<15> dmem_addr<16> dmem_addr<15> rd_mux_sel<1> rd_mux_sel<2> rd_sel<31> rs1_sel<31> rs2_sel<31> rd_sel<30> rs1_sel<30>
+ rs2_sel<30> rd_sel<29> rs1_sel<29> rs2_sel<29> rd_sel<28> rs1_sel<28> rs2_sel<28> rd_sel<27> rs1_sel<27> rs2_sel<27> rd_sel<26> rs1_sel<26> rs2_sel<26> rd_sel<25> rs1_sel<25> rs2_sel<25> rd_sel<24> rs1_sel<24> rs2_sel<24> rd_sel<23>
+ rs1_sel<23> rs2_sel<23> rd_sel<22> rs1_sel<22> rs2_sel<22> rd_sel<21> rs1_sel<21> rs2_sel<21> rd_sel<20> rs1_sel<20> rs2_sel<20> rd_sel<19> rs1_sel<19> rs2_sel<19> rd_sel<18> rs1_sel<18> rs2_sel<18> rd_sel<17> rs1_sel<17> rs2_sel<17>
+ rd_sel<16> rs1_sel<16> rs2_sel<16> rd_sel<15> rs1_sel<15> rs2_sel<15> rd_sel<14> rs1_sel<14> rs2_sel<14> rd_sel<13> rs1_sel<13> rs2_sel<13> rd_sel<12> rs1_sel<12> rs2_sel<12> rd_sel<11> rs1_sel<11> rs2_sel<11> rd_sel<10> rs1_sel<10>
+ rs2_sel<10> rd_sel<9> rs1_sel<9> rs2_sel<9> rd_sel<8> rs1_sel<8> rs2_sel<8> rd_sel<7> rs1_sel<7> rs2_sel<7> rd_sel<6> rs1_sel<6> rs2_sel<6> rd_sel<5> rs1_sel<5> rs2_sel<5> rd_sel<4> rs1_sel<4> rs2_sel<4> rd_sel<3>
+ rs1_sel<3> rs2_sel<3> rd_sel<2> rs1_sel<2> rs2_sel<2> rd_sel<1> rs1_sel<1> 235 rs2_sel<1> rs2_sel<0> rs1_sel<0> clk 244 336 338 dmem_wdata<16> dmem_wdata<15> 286 288 alu_mux_1_sel
+ imem_addr<16> imem_addr<15> alu_inv_rs2 alu_mux_2_sel 316 342 234 alu_op<0> alu_op<1> shift_dir 321 320 348 346 296 291 349 343 237 147
+ 6 337 339 164 shift_msb 351 146 148 322 317 149 153 157 354 158 cmp_mux_sel 350 323 352 326
+ 327 353 pc_mux_sel rst
+ ICV_31 $T=0 0 0 0 $X=0 $Y=67600
X8 mem_mux_sel<0> dmem_rdata<20> dmem_rdata<19> dmem_rdata<18> dmem_rdata<17> dmem_rdata<7> dmem_rdata<15> vss! mem_mux_sel<1> mem_mux_sel<2> vdd! rd_mux_sel<0> imm<20> imm<19> imm<18> imm<17> dmem_addr<20> dmem_addr<19> dmem_addr<18> dmem_addr<17>
+ rd_mux_sel<1> rd_mux_sel<2> rd_sel<31> rs1_sel<31> rs2_sel<31> rd_sel<30> rs1_sel<30> rs2_sel<30> rd_sel<29> rs1_sel<29> rs2_sel<29> rd_sel<28> rs1_sel<28> rs2_sel<28> rd_sel<27> rs1_sel<27> rs2_sel<27> rd_sel<26> rs1_sel<26> rs2_sel<26>
+ rd_sel<25> rs1_sel<25> rs2_sel<25> rd_sel<24> rs1_sel<24> rs2_sel<24> rd_sel<23> rs1_sel<23> rs2_sel<23> rd_sel<22> rs1_sel<22> rs2_sel<22> rd_sel<21> rs1_sel<21> rs2_sel<21> rd_sel<20> rs1_sel<20> rs2_sel<20> rd_sel<19> rs1_sel<19>
+ rs2_sel<19> rd_sel<18> rs1_sel<18> rs2_sel<18> rd_sel<17> rs1_sel<17> rs2_sel<17> rd_sel<16> rs1_sel<16> rs2_sel<16> rd_sel<15> rs1_sel<15> rs2_sel<15> rd_sel<14> rs1_sel<14> rs2_sel<14> rd_sel<13> rs1_sel<13> rs2_sel<13> rd_sel<12>
+ rs1_sel<12> rs2_sel<12> rd_sel<11> rs1_sel<11> rs2_sel<11> rd_sel<10> rs1_sel<10> rs2_sel<10> rd_sel<9> rs1_sel<9> rs2_sel<9> rd_sel<8> rs1_sel<8> rs2_sel<8> rd_sel<7> rs1_sel<7> rs2_sel<7> rd_sel<6> rs1_sel<6> rs2_sel<6>
+ rd_sel<5> rs1_sel<5> rs2_sel<5> rd_sel<4> rs1_sel<4> rs2_sel<4> rd_sel<3> rs1_sel<3> rs2_sel<3> rd_sel<2> rs1_sel<2> 289 260 rs2_sel<2> rd_sel<1> rs1_sel<1> 262 365 367 rs2_sel<1>
+ rs2_sel<0> rs1_sel<0> 369 clk 338 310 312 dmem_wdata<20> dmem_wdata<19> dmem_wdata<18> dmem_wdata<17> alu_mux_1_sel imem_addr<20> imem_addr<19> imem_addr<18> imem_addr<17> alu_inv_rs2 alu_mux_2_sel 342 375
+ 286 261 288 alu_op<0> alu_op<1> shift_dir 348 346 382 386 349 343 322 317 383 377 387 376 263 384
+ 193 192 163 7 385 366 368 370 199 198 167 8 shift_msb 146 149 336 153 287 157 194
+ 190 154 155 158 cmp_mux_sel 388 350 389 352 353 390 pc_mux_sel rst
+ ICV_36 $T=0 0 0 0 $X=0 $Y=50930
X9 mem_mux_sel<0> dmem_rdata<22> dmem_rdata<21> dmem_rdata<7> dmem_rdata<15> vss! mem_mux_sel<1> mem_mux_sel<2> vdd! rd_mux_sel<0> imm<22> imm<21> dmem_addr<22> dmem_addr<21> rd_mux_sel<1> rd_mux_sel<2> rd_sel<31> rs1_sel<31> rs2_sel<31> rd_sel<30>
+ rs1_sel<30> rs2_sel<30> rd_sel<29> rs1_sel<29> rs2_sel<29> rd_sel<28> rs1_sel<28> rs2_sel<28> rd_sel<27> rs1_sel<27> rs2_sel<27> rd_sel<26> rs1_sel<26> rs2_sel<26> rd_sel<25> rs1_sel<25> rs2_sel<25> rd_sel<24> rs1_sel<24> rs2_sel<24>
+ rd_sel<23> rs1_sel<23> rs2_sel<23> rd_sel<22> rs1_sel<22> rs2_sel<22> rd_sel<21> rs1_sel<21> rs2_sel<21> rd_sel<20> rs1_sel<20> rs2_sel<20> rd_sel<19> rs1_sel<19> rs2_sel<19> rd_sel<18> rs1_sel<18> rs2_sel<18> rd_sel<17> rs1_sel<17>
+ rs2_sel<17> rd_sel<16> rs1_sel<16> rs2_sel<16> rd_sel<15> rs1_sel<15> rs2_sel<15> rd_sel<14> rs1_sel<14> rs2_sel<14> rd_sel<13> rs1_sel<13> rs2_sel<13> rd_sel<12> rs1_sel<12> rs2_sel<12> rd_sel<11> rs1_sel<11> rs2_sel<11> rd_sel<10>
+ rs1_sel<10> rs2_sel<10> rd_sel<9> rs1_sel<9> rs2_sel<9> rd_sel<8> rs1_sel<8> rs2_sel<8> rd_sel<7> rs1_sel<7> rs2_sel<7> rd_sel<6> rs1_sel<6> rs2_sel<6> rd_sel<5> rs1_sel<5> rs2_sel<5> rd_sel<4> rs1_sel<4> rs2_sel<4>
+ rd_sel<3> rs1_sel<3> rs2_sel<3> rd_sel<2> rs1_sel<2> 313 399 rs2_sel<2> rd_sel<1> rs1_sel<1> rs2_sel<1> rs2_sel<0> rs1_sel<0> 369 clk dmem_wdata<22> dmem_wdata<21> alu_mux_1_sel imem_addr<22> imem_addr<21>
+ alu_inv_rs2 alu_mux_2_sel 375 403 312 310 alu_op<0> alu_op<1> shift_dir 382 386 407 411 387 376 408 404 409 220 217
+ 410 400 224 225 shift_msb 146 383 377 149 367 153 311 157 9 218 158 cmp_mux_sel 10 388 11
+ 389 390 412 pc_mux_sel rst
+ ICV_37 $T=0 0 0 0 $X=0 $Y=41600
X10 mem_mux_sel<0> dmem_rdata<24> dmem_rdata<23> dmem_rdata<7> dmem_rdata<15> vss! mem_mux_sel<1> mem_mux_sel<2> vdd! rd_mux_sel<0> imm<24> imm<23> dmem_addr<24> dmem_addr<23> rd_mux_sel<1> rd_mux_sel<2> rd_sel<31> rs1_sel<31> rs2_sel<31> rd_sel<30>
+ rs1_sel<30> rs2_sel<30> rd_sel<29> rs1_sel<29> rs2_sel<29> rd_sel<28> rs1_sel<28> rs2_sel<28> rd_sel<27> rs1_sel<27> rs2_sel<27> rd_sel<26> rs1_sel<26> rs2_sel<26> rd_sel<25> rs1_sel<25> rs2_sel<25> rd_sel<24> rs1_sel<24> rs2_sel<24>
+ rd_sel<23> rs1_sel<23> rs2_sel<23> rd_sel<22> rs1_sel<22> rs2_sel<22> rd_sel<21> rs1_sel<21> rs2_sel<21> rd_sel<20> rs1_sel<20> rs2_sel<20> rd_sel<19> rs1_sel<19> rs2_sel<19> rd_sel<18> rs1_sel<18> rs2_sel<18> rd_sel<17> rs1_sel<17>
+ rs2_sel<17> rd_sel<16> rs1_sel<16> rs2_sel<16> rd_sel<15> rs1_sel<15> rs2_sel<15> rd_sel<14> rs1_sel<14> rs2_sel<14> rd_sel<13> rs1_sel<13> rs2_sel<13> rd_sel<12> rs1_sel<12> rs2_sel<12> rd_sel<11> rs1_sel<11> rs2_sel<11> rd_sel<10>
+ rs1_sel<10> rs2_sel<10> rd_sel<9> rs1_sel<9> rs2_sel<9> rd_sel<8> rs1_sel<8> rs2_sel<8> rd_sel<7> rs1_sel<7> rs2_sel<7> rd_sel<6> rs1_sel<6> rs2_sel<6> rd_sel<5> rs1_sel<5> rs2_sel<5> rd_sel<4> rs1_sel<4> rs2_sel<4>
+ rd_sel<3> rs1_sel<3> rs2_sel<3> rd_sel<2> rs1_sel<2> 339 419 rs2_sel<2> rd_sel<1> rs1_sel<1> 365 rs2_sel<1> rs2_sel<0> rs1_sel<0> clk dmem_wdata<24> dmem_wdata<23> alu_mux_1_sel imem_addr<24> imem_addr<23>
+ alu_inv_rs2 alu_mux_2_sel 403 423 336 338 alu_op<0> alu_op<1> shift_dir 407 411 427 430 383 377 428 424 429 235 244
+ shift_msb 420 250 251 146 408 404 149 384 153 337 157 247 246 158 cmp_mux_sel 431 10 12 11
+ 412 432 pc_mux_sel rst
+ ICV_38 $T=0 0 0 0 $X=0 $Y=32400
X11 mem_mux_sel<0> dmem_rdata<26> dmem_rdata<25> dmem_rdata<7> dmem_rdata<15> vss! mem_mux_sel<1> mem_mux_sel<2> vdd! rd_mux_sel<0> imm<26> imm<25> dmem_addr<26> dmem_addr<25> rd_mux_sel<1> rd_mux_sel<2> rd_sel<31> rs1_sel<31> rs2_sel<31> rd_sel<30>
+ rs1_sel<30> rs2_sel<30> rd_sel<29> rs1_sel<29> rs2_sel<29> rd_sel<28> rs1_sel<28> rs2_sel<28> rd_sel<27> rs1_sel<27> rs2_sel<27> rd_sel<26> rs1_sel<26> rs2_sel<26> rd_sel<25> rs1_sel<25> rs2_sel<25> rd_sel<24> rs1_sel<24> rs2_sel<24>
+ rd_sel<23> rs1_sel<23> rs2_sel<23> rd_sel<22> rs1_sel<22> rs2_sel<22> rd_sel<21> rs1_sel<21> rs2_sel<21> rd_sel<20> rs1_sel<20> rs2_sel<20> rd_sel<19> rs1_sel<19> rs2_sel<19> rd_sel<18> rs1_sel<18> rs2_sel<18> rd_sel<17> rs1_sel<17>
+ rs2_sel<17> rd_sel<16> rs1_sel<16> rs2_sel<16> rd_sel<15> rs1_sel<15> rs2_sel<15> rd_sel<14> rs1_sel<14> rs2_sel<14> rd_sel<13> rs1_sel<13> rs2_sel<13> rd_sel<12> rs1_sel<12> rs2_sel<12> rd_sel<11> rs1_sel<11> rs2_sel<11> rd_sel<10>
+ rs1_sel<10> rs2_sel<10> rd_sel<9> rs1_sel<9> rs2_sel<9> rd_sel<8> rs1_sel<8> rs2_sel<8> rd_sel<7> rs1_sel<7> rs2_sel<7> rd_sel<6> rs1_sel<6> rs2_sel<6> rd_sel<5> rs1_sel<5> rs2_sel<5> rd_sel<4> rs1_sel<4> rs2_sel<4>
+ rd_sel<3> rs1_sel<3> rs2_sel<3> rd_sel<2> rs1_sel<2> 399 rs2_sel<2> rd_sel<1> rs1_sel<1> rs2_sel<1> rs2_sel<0> rs1_sel<0> 370 clk dmem_wdata<26> dmem_wdata<25> alu_mux_1_sel imem_addr<26> imem_addr<25> alu_inv_rs2
+ alu_mux_2_sel 423 441 369 367 alu_op<0> alu_op<1> shift_dir 427 430 445 448 408 404 446 442 447 449 260 262
+ shift_msb 277 276 146 428 424 149 409 153 368 157 273 272 158 cmp_mux_sel 450 431 451 12 432
+ 452 pc_mux_sel rst
+ ICV_39 $T=0 0 0 0 $X=0 $Y=23150
X12 mem_mux_sel<0> dmem_rdata<28> dmem_rdata<27> dmem_rdata<7> dmem_rdata<15> vss! mem_mux_sel<1> mem_mux_sel<2> vdd! rd_mux_sel<0> imm<28> imm<27> dmem_addr<28> dmem_addr<27> rd_mux_sel<1> rd_mux_sel<2> rd_sel<31> rs1_sel<31> rs2_sel<31> rd_sel<30>
+ rs1_sel<30> rs2_sel<30> rd_sel<29> rs1_sel<29> rs2_sel<29> rd_sel<28> rs1_sel<28> rs2_sel<28> rd_sel<27> rs1_sel<27> rs2_sel<27> rd_sel<26> rs1_sel<26> rs2_sel<26> rd_sel<25> rs1_sel<25> rs2_sel<25> rd_sel<24> rs1_sel<24> rs2_sel<24>
+ rd_sel<23> rs1_sel<23> rs2_sel<23> rd_sel<22> rs1_sel<22> rs2_sel<22> rd_sel<21> rs1_sel<21> rs2_sel<21> rd_sel<20> rs1_sel<20> rs2_sel<20> rd_sel<19> rs1_sel<19> rs2_sel<19> rd_sel<18> rs1_sel<18> rs2_sel<18> rd_sel<17> rs1_sel<17>
+ rs2_sel<17> rd_sel<16> rs1_sel<16> rs2_sel<16> rd_sel<15> rs1_sel<15> rs2_sel<15> rd_sel<14> rs1_sel<14> rs2_sel<14> rd_sel<13> rs1_sel<13> rs2_sel<13> rd_sel<12> rs1_sel<12> rs2_sel<12> rd_sel<11> rs1_sel<11> rs2_sel<11> rd_sel<10>
+ rs1_sel<10> rs2_sel<10> rd_sel<9> rs1_sel<9> rs2_sel<9> rd_sel<8> rs1_sel<8> rs2_sel<8> rd_sel<7> rs1_sel<7> rs2_sel<7> rd_sel<6> rs1_sel<6> rs2_sel<6> rd_sel<5> rs1_sel<5> rs2_sel<5> rd_sel<4> rs1_sel<4> rs2_sel<4>
+ rd_sel<3> rs1_sel<3> rs2_sel<3> rd_sel<2> rs1_sel<2> 419 rs2_sel<2> rd_sel<1> rs1_sel<1> 366 rs2_sel<1> rs2_sel<0> rs1_sel<0> clk dmem_wdata<28> dmem_wdata<27> alu_mux_1_sel imem_addr<28> imem_addr<27> alu_inv_rs2
+ alu_mux_2_sel 441 461 384 365 alu_op<0> alu_op<1> shift_dir 445 448 465 467 428 424 466 462 shift_msb 468 287 289
+ 303 302 146 446 442 149 429 153 385 157 299 298 158 cmp_mux_sel 469 450 13 451 452 470
+ pc_mux_sel rst
+ ICV_40 $T=0 0 0 0 $X=0 $Y=13800
X13 mem_mux_sel<0> dmem_rdata<31> dmem_rdata<30> dmem_rdata<29> dmem_rdata<7> dmem_rdata<15> vss! mem_mux_sel<1> mem_mux_sel<2> vdd! rd_mux_sel<0> imm<31> imm<30> imm<29> dmem_addr<31> dmem_addr<30> dmem_addr<29> rd_mux_sel<1> rd_mux_sel<2> rd_sel<31>
+ rs1_sel<31> rs2_sel<31> rd_sel<30> rs1_sel<30> rs2_sel<30> rd_sel<29> rs1_sel<29> rs2_sel<29> rd_sel<28> rs1_sel<28> rs2_sel<28> rd_sel<27> rs1_sel<27> rs2_sel<27> rd_sel<26> rs1_sel<26> rs2_sel<26> rd_sel<25> rs1_sel<25> rs2_sel<25>
+ rd_sel<24> rs1_sel<24> rs2_sel<24> rd_sel<23> rs1_sel<23> rs2_sel<23> rd_sel<22> rs1_sel<22> rs2_sel<22> rd_sel<21> rs1_sel<21> rs2_sel<21> rd_sel<20> rs1_sel<20> rs2_sel<20> rd_sel<19> rs1_sel<19> rs2_sel<19> rd_sel<18> rs1_sel<18>
+ rs2_sel<18> rd_sel<17> rs1_sel<17> rs2_sel<17> rd_sel<16> rs1_sel<16> rs2_sel<16> rd_sel<15> rs1_sel<15> rs2_sel<15> rd_sel<14> rs1_sel<14> rs2_sel<14> rd_sel<13> rs1_sel<13> rs2_sel<13> rd_sel<12> rs1_sel<12> rs2_sel<12> rd_sel<11>
+ rs1_sel<11> rs2_sel<11> rd_sel<10> rs1_sel<10> rs2_sel<10> rd_sel<9> rs1_sel<9> rs2_sel<9> rd_sel<8> rs1_sel<8> rs2_sel<8> rd_sel<7> rs1_sel<7> rs2_sel<7> rd_sel<6> rs1_sel<6> rs2_sel<6> rd_sel<5> rs1_sel<5> rs2_sel<5>
+ rd_sel<4> rs1_sel<4> rs2_sel<4> rd_sel<3> rs1_sel<3> rs2_sel<3> rd_sel<2> rs1_sel<2> 400 420 rs2_sel<2> rd_sel<1> rs1_sel<1> 410 rs2_sel<1> rs2_sel<0> rs1_sel<0> clk cmp_a_31 dmem_wdata<31>
+ dmem_wdata<30> dmem_wdata<29> alu_mux_1_sel imem_addr<31> imem_addr<30> imem_addr<29> alu_inv_rs2 alu_mux_2_sel 461 399 409 419 alu_op<0> alu_op<1> shift_dir 465 467 shift_msb 462 446
+ 442 339 311 313 354 329 328 146 466 149 468 447 449 153 157 351 325 324 158 cmp_mux_sel
+ cmp_b_31 469 13 470 pc_mux_sel rst
+ ICV_41 $T=0 0 0 0 $X=0 $Y=0
.ENDS
***************************************
