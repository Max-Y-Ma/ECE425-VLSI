* SPICE NETLIST
***************************************

.SUBCKT M1_POLY_CDNS_711421196622
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NTAP_CDNS_711421196621
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT PTAP_CDNS_711421196620
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_1
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_2
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_3
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_4
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_5
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_6
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_7
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_8
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_9
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_10
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_11
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_12
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_13
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_14
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_15
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_16
** N=1 EP=0 IP=3 FDC=0
.ENDS
***************************************
.SUBCKT ICV_17
** N=1 EP=0 IP=3 FDC=0
.ENDS
***************************************
.SUBCKT ICV_18
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_19
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_20
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_21
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_22
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_23
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_24 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168
** N=1109 EP=168 IP=2241 FDC=2700
M0 170 1 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=134870 $D=1
M1 171 1 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=139500 $D=1
M2 172 1 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=144130 $D=1
M3 173 170 2 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=134870 $D=1
M4 174 171 3 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=139500 $D=1
M5 175 172 4 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=144130 $D=1
M6 8 1 173 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=134870 $D=1
M7 9 1 174 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=139500 $D=1
M8 136 1 175 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=144130 $D=1
M9 176 170 2 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=134870 $D=1
M10 177 171 3 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=139500 $D=1
M11 178 172 4 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=144130 $D=1
M12 2 1 176 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=134870 $D=1
M13 3 1 177 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=139500 $D=1
M14 4 1 178 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=144130 $D=1
M15 179 170 2 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=134870 $D=1
M16 180 171 3 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=139500 $D=1
M17 181 172 4 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=144130 $D=1
M18 2 1 179 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=134870 $D=1
M19 3 1 180 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=139500 $D=1
M20 4 1 181 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=144130 $D=1
M21 185 182 179 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=134870 $D=1
M22 186 183 180 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=139500 $D=1
M23 187 184 181 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=144130 $D=1
M24 182 5 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=134870 $D=1
M25 183 5 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=139500 $D=1
M26 184 5 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=144130 $D=1
M27 188 182 176 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=134870 $D=1
M28 189 183 177 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=139500 $D=1
M29 190 184 178 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=144130 $D=1
M30 173 5 188 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=134870 $D=1
M31 174 5 189 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=139500 $D=1
M32 175 5 190 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=144130 $D=1
M33 191 6 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=134870 $D=1
M34 192 6 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=139500 $D=1
M35 193 6 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=144130 $D=1
M36 194 191 188 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=134870 $D=1
M37 195 192 189 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=139500 $D=1
M38 196 193 190 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=144130 $D=1
M39 185 6 194 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=134870 $D=1
M40 186 6 195 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=139500 $D=1
M41 187 6 196 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=144130 $D=1
M42 197 7 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=134870 $D=1
M43 198 7 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=139500 $D=1
M44 199 7 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=144130 $D=1
M45 200 197 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=134870 $D=1
M46 201 198 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=139500 $D=1
M47 202 199 10 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=144130 $D=1
M48 11 7 200 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=134870 $D=1
M49 12 7 201 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=139500 $D=1
M50 13 7 202 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=144130 $D=1
M51 203 197 14 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=134870 $D=1
M52 204 198 15 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=139500 $D=1
M53 205 199 16 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=144130 $D=1
M54 206 7 203 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=134870 $D=1
M55 207 7 204 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=139500 $D=1
M56 208 7 205 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=144130 $D=1
M57 212 197 209 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=134870 $D=1
M58 213 198 210 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=139500 $D=1
M59 214 199 211 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=144130 $D=1
M60 194 7 212 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=134870 $D=1
M61 195 7 213 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=139500 $D=1
M62 196 7 214 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=144130 $D=1
M63 218 215 212 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=134870 $D=1
M64 219 216 213 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=139500 $D=1
M65 220 217 214 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=144130 $D=1
M66 215 17 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=134870 $D=1
M67 216 17 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=139500 $D=1
M68 217 17 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=144130 $D=1
M69 221 215 203 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=134870 $D=1
M70 222 216 204 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=139500 $D=1
M71 223 217 205 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=144130 $D=1
M72 200 17 221 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=134870 $D=1
M73 201 17 222 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=139500 $D=1
M74 202 17 223 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=144130 $D=1
M75 224 18 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=134870 $D=1
M76 225 18 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=139500 $D=1
M77 226 18 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=144130 $D=1
M78 227 224 221 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=134870 $D=1
M79 228 225 222 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=139500 $D=1
M80 229 226 223 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=144130 $D=1
M81 218 18 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=134870 $D=1
M82 219 18 228 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=139500 $D=1
M83 220 18 229 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=144130 $D=1
M84 8 19 230 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=134870 $D=1
M85 9 19 231 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=139500 $D=1
M86 136 19 232 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=144130 $D=1
M87 233 20 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=134870 $D=1
M88 234 20 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=139500 $D=1
M89 235 20 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=144130 $D=1
M90 236 19 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=134870 $D=1
M91 237 19 228 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=139500 $D=1
M92 238 19 229 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=144130 $D=1
M93 8 236 945 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=134870 $D=1
M94 9 237 946 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=139500 $D=1
M95 136 238 947 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=144130 $D=1
M96 239 945 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=134870 $D=1
M97 240 946 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=139500 $D=1
M98 241 947 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=144130 $D=1
M99 236 230 239 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=134870 $D=1
M100 237 231 240 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=139500 $D=1
M101 238 232 241 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=144130 $D=1
M102 239 20 242 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=134870 $D=1
M103 240 20 243 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=139500 $D=1
M104 241 20 244 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=144130 $D=1
M105 248 21 239 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=134870 $D=1
M106 249 21 240 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=139500 $D=1
M107 250 21 241 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=144130 $D=1
M108 245 21 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=134870 $D=1
M109 246 21 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=139500 $D=1
M110 247 21 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=144130 $D=1
M111 8 22 251 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=134870 $D=1
M112 9 22 252 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=139500 $D=1
M113 136 22 253 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=144130 $D=1
M114 254 23 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=134870 $D=1
M115 255 23 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=139500 $D=1
M116 256 23 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=144130 $D=1
M117 257 22 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=134870 $D=1
M118 258 22 228 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=139500 $D=1
M119 259 22 229 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=144130 $D=1
M120 8 257 948 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=134870 $D=1
M121 9 258 949 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=139500 $D=1
M122 136 259 950 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=144130 $D=1
M123 260 948 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=134870 $D=1
M124 261 949 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=139500 $D=1
M125 262 950 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=144130 $D=1
M126 257 251 260 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=134870 $D=1
M127 258 252 261 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=139500 $D=1
M128 259 253 262 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=144130 $D=1
M129 260 23 242 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=134870 $D=1
M130 261 23 243 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=139500 $D=1
M131 262 23 244 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=144130 $D=1
M132 248 24 260 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=134870 $D=1
M133 249 24 261 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=139500 $D=1
M134 250 24 262 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=144130 $D=1
M135 263 24 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=134870 $D=1
M136 264 24 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=139500 $D=1
M137 265 24 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=144130 $D=1
M138 8 25 266 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=134870 $D=1
M139 9 25 267 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=139500 $D=1
M140 136 25 268 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=144130 $D=1
M141 269 26 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=134870 $D=1
M142 270 26 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=139500 $D=1
M143 271 26 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=144130 $D=1
M144 272 25 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=134870 $D=1
M145 273 25 228 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=139500 $D=1
M146 274 25 229 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=144130 $D=1
M147 8 272 951 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=134870 $D=1
M148 9 273 952 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=139500 $D=1
M149 136 274 953 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=144130 $D=1
M150 275 951 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=134870 $D=1
M151 276 952 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=139500 $D=1
M152 277 953 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=144130 $D=1
M153 272 266 275 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=134870 $D=1
M154 273 267 276 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=139500 $D=1
M155 274 268 277 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=144130 $D=1
M156 275 26 242 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=134870 $D=1
M157 276 26 243 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=139500 $D=1
M158 277 26 244 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=144130 $D=1
M159 248 27 275 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=134870 $D=1
M160 249 27 276 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=139500 $D=1
M161 250 27 277 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=144130 $D=1
M162 278 27 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=134870 $D=1
M163 279 27 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=139500 $D=1
M164 280 27 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=144130 $D=1
M165 8 28 281 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=134870 $D=1
M166 9 28 282 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=139500 $D=1
M167 136 28 283 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=144130 $D=1
M168 284 29 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=134870 $D=1
M169 285 29 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=139500 $D=1
M170 286 29 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=144130 $D=1
M171 287 28 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=134870 $D=1
M172 288 28 228 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=139500 $D=1
M173 289 28 229 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=144130 $D=1
M174 8 287 954 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=134870 $D=1
M175 9 288 955 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=139500 $D=1
M176 136 289 956 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=144130 $D=1
M177 290 954 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=134870 $D=1
M178 291 955 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=139500 $D=1
M179 292 956 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=144130 $D=1
M180 287 281 290 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=134870 $D=1
M181 288 282 291 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=139500 $D=1
M182 289 283 292 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=144130 $D=1
M183 290 29 242 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=134870 $D=1
M184 291 29 243 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=139500 $D=1
M185 292 29 244 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=144130 $D=1
M186 248 30 290 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=134870 $D=1
M187 249 30 291 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=139500 $D=1
M188 250 30 292 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=144130 $D=1
M189 293 30 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=134870 $D=1
M190 294 30 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=139500 $D=1
M191 295 30 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=144130 $D=1
M192 8 31 296 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=134870 $D=1
M193 9 31 297 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=139500 $D=1
M194 136 31 298 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=144130 $D=1
M195 299 32 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=134870 $D=1
M196 300 32 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=139500 $D=1
M197 301 32 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=144130 $D=1
M198 302 31 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=134870 $D=1
M199 303 31 228 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=139500 $D=1
M200 304 31 229 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=144130 $D=1
M201 8 302 957 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=134870 $D=1
M202 9 303 958 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=139500 $D=1
M203 136 304 959 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=144130 $D=1
M204 305 957 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=134870 $D=1
M205 306 958 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=139500 $D=1
M206 307 959 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=144130 $D=1
M207 302 296 305 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=134870 $D=1
M208 303 297 306 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=139500 $D=1
M209 304 298 307 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=144130 $D=1
M210 305 32 242 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=134870 $D=1
M211 306 32 243 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=139500 $D=1
M212 307 32 244 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=144130 $D=1
M213 248 33 305 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=134870 $D=1
M214 249 33 306 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=139500 $D=1
M215 250 33 307 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=144130 $D=1
M216 308 33 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=134870 $D=1
M217 309 33 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=139500 $D=1
M218 310 33 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=144130 $D=1
M219 8 34 311 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=134870 $D=1
M220 9 34 312 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=139500 $D=1
M221 136 34 313 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=144130 $D=1
M222 314 35 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=134870 $D=1
M223 315 35 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=139500 $D=1
M224 316 35 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=144130 $D=1
M225 317 34 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=134870 $D=1
M226 318 34 228 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=139500 $D=1
M227 319 34 229 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=144130 $D=1
M228 8 317 960 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=134870 $D=1
M229 9 318 961 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=139500 $D=1
M230 136 319 962 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=144130 $D=1
M231 320 960 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=134870 $D=1
M232 321 961 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=139500 $D=1
M233 322 962 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=144130 $D=1
M234 317 311 320 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=134870 $D=1
M235 318 312 321 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=139500 $D=1
M236 319 313 322 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=144130 $D=1
M237 320 35 242 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=134870 $D=1
M238 321 35 243 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=139500 $D=1
M239 322 35 244 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=144130 $D=1
M240 248 36 320 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=134870 $D=1
M241 249 36 321 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=139500 $D=1
M242 250 36 322 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=144130 $D=1
M243 323 36 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=134870 $D=1
M244 324 36 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=139500 $D=1
M245 325 36 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=144130 $D=1
M246 8 37 326 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=134870 $D=1
M247 9 37 327 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=139500 $D=1
M248 136 37 328 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=144130 $D=1
M249 329 38 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=134870 $D=1
M250 330 38 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=139500 $D=1
M251 331 38 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=144130 $D=1
M252 332 37 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=134870 $D=1
M253 333 37 228 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=139500 $D=1
M254 334 37 229 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=144130 $D=1
M255 8 332 963 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=134870 $D=1
M256 9 333 964 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=139500 $D=1
M257 136 334 965 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=144130 $D=1
M258 335 963 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=134870 $D=1
M259 336 964 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=139500 $D=1
M260 337 965 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=144130 $D=1
M261 332 326 335 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=134870 $D=1
M262 333 327 336 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=139500 $D=1
M263 334 328 337 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=144130 $D=1
M264 335 38 242 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=134870 $D=1
M265 336 38 243 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=139500 $D=1
M266 337 38 244 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=144130 $D=1
M267 248 39 335 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=134870 $D=1
M268 249 39 336 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=139500 $D=1
M269 250 39 337 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=144130 $D=1
M270 338 39 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=134870 $D=1
M271 339 39 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=139500 $D=1
M272 340 39 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=144130 $D=1
M273 8 40 341 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=134870 $D=1
M274 9 40 342 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=139500 $D=1
M275 136 40 343 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=144130 $D=1
M276 344 41 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=134870 $D=1
M277 345 41 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=139500 $D=1
M278 346 41 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=144130 $D=1
M279 347 40 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=134870 $D=1
M280 348 40 228 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=139500 $D=1
M281 349 40 229 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=144130 $D=1
M282 8 347 966 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=134870 $D=1
M283 9 348 967 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=139500 $D=1
M284 136 349 968 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=144130 $D=1
M285 350 966 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=134870 $D=1
M286 351 967 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=139500 $D=1
M287 352 968 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=144130 $D=1
M288 347 341 350 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=134870 $D=1
M289 348 342 351 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=139500 $D=1
M290 349 343 352 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=144130 $D=1
M291 350 41 242 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=134870 $D=1
M292 351 41 243 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=139500 $D=1
M293 352 41 244 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=144130 $D=1
M294 248 42 350 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=134870 $D=1
M295 249 42 351 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=139500 $D=1
M296 250 42 352 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=144130 $D=1
M297 353 42 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=134870 $D=1
M298 354 42 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=139500 $D=1
M299 355 42 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=144130 $D=1
M300 8 43 356 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=134870 $D=1
M301 9 43 357 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=139500 $D=1
M302 136 43 358 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=144130 $D=1
M303 359 44 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=134870 $D=1
M304 360 44 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=139500 $D=1
M305 361 44 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=144130 $D=1
M306 362 43 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=134870 $D=1
M307 363 43 228 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=139500 $D=1
M308 364 43 229 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=144130 $D=1
M309 8 362 969 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=134870 $D=1
M310 9 363 970 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=139500 $D=1
M311 136 364 971 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=144130 $D=1
M312 365 969 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=134870 $D=1
M313 366 970 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=139500 $D=1
M314 367 971 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=144130 $D=1
M315 362 356 365 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=134870 $D=1
M316 363 357 366 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=139500 $D=1
M317 364 358 367 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=144130 $D=1
M318 365 44 242 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=134870 $D=1
M319 366 44 243 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=139500 $D=1
M320 367 44 244 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=144130 $D=1
M321 248 45 365 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=134870 $D=1
M322 249 45 366 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=139500 $D=1
M323 250 45 367 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=144130 $D=1
M324 368 45 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=134870 $D=1
M325 369 45 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=139500 $D=1
M326 370 45 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=144130 $D=1
M327 8 46 371 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=134870 $D=1
M328 9 46 372 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=139500 $D=1
M329 136 46 373 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=144130 $D=1
M330 374 47 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=134870 $D=1
M331 375 47 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=139500 $D=1
M332 376 47 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=144130 $D=1
M333 377 46 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=134870 $D=1
M334 378 46 228 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=139500 $D=1
M335 379 46 229 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=144130 $D=1
M336 8 377 972 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=134870 $D=1
M337 9 378 973 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=139500 $D=1
M338 136 379 974 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=144130 $D=1
M339 380 972 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=134870 $D=1
M340 381 973 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=139500 $D=1
M341 382 974 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=144130 $D=1
M342 377 371 380 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=134870 $D=1
M343 378 372 381 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=139500 $D=1
M344 379 373 382 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=144130 $D=1
M345 380 47 242 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=134870 $D=1
M346 381 47 243 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=139500 $D=1
M347 382 47 244 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=144130 $D=1
M348 248 48 380 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=134870 $D=1
M349 249 48 381 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=139500 $D=1
M350 250 48 382 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=144130 $D=1
M351 383 48 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=134870 $D=1
M352 384 48 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=139500 $D=1
M353 385 48 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=144130 $D=1
M354 8 49 386 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=134870 $D=1
M355 9 49 387 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=139500 $D=1
M356 136 49 388 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=144130 $D=1
M357 389 50 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=134870 $D=1
M358 390 50 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=139500 $D=1
M359 391 50 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=144130 $D=1
M360 392 49 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=134870 $D=1
M361 393 49 228 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=139500 $D=1
M362 394 49 229 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=144130 $D=1
M363 8 392 975 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=134870 $D=1
M364 9 393 976 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=139500 $D=1
M365 136 394 977 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=144130 $D=1
M366 395 975 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=134870 $D=1
M367 396 976 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=139500 $D=1
M368 397 977 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=144130 $D=1
M369 392 386 395 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=134870 $D=1
M370 393 387 396 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=139500 $D=1
M371 394 388 397 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=144130 $D=1
M372 395 50 242 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=134870 $D=1
M373 396 50 243 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=139500 $D=1
M374 397 50 244 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=144130 $D=1
M375 248 51 395 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=134870 $D=1
M376 249 51 396 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=139500 $D=1
M377 250 51 397 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=144130 $D=1
M378 398 51 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=134870 $D=1
M379 399 51 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=139500 $D=1
M380 400 51 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=144130 $D=1
M381 8 52 401 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=134870 $D=1
M382 9 52 402 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=139500 $D=1
M383 136 52 403 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=144130 $D=1
M384 404 53 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=134870 $D=1
M385 405 53 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=139500 $D=1
M386 406 53 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=144130 $D=1
M387 407 52 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=134870 $D=1
M388 408 52 228 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=139500 $D=1
M389 409 52 229 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=144130 $D=1
M390 8 407 978 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=134870 $D=1
M391 9 408 979 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=139500 $D=1
M392 136 409 980 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=144130 $D=1
M393 410 978 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=134870 $D=1
M394 411 979 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=139500 $D=1
M395 412 980 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=144130 $D=1
M396 407 401 410 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=134870 $D=1
M397 408 402 411 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=139500 $D=1
M398 409 403 412 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=144130 $D=1
M399 410 53 242 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=134870 $D=1
M400 411 53 243 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=139500 $D=1
M401 412 53 244 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=144130 $D=1
M402 248 54 410 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=134870 $D=1
M403 249 54 411 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=139500 $D=1
M404 250 54 412 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=144130 $D=1
M405 413 54 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=134870 $D=1
M406 414 54 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=139500 $D=1
M407 415 54 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=144130 $D=1
M408 8 55 416 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=134870 $D=1
M409 9 55 417 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=139500 $D=1
M410 136 55 418 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=144130 $D=1
M411 419 56 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=134870 $D=1
M412 420 56 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=139500 $D=1
M413 421 56 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=144130 $D=1
M414 422 55 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=134870 $D=1
M415 423 55 228 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=139500 $D=1
M416 424 55 229 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=144130 $D=1
M417 8 422 981 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=134870 $D=1
M418 9 423 982 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=139500 $D=1
M419 136 424 983 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=144130 $D=1
M420 425 981 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=134870 $D=1
M421 426 982 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=139500 $D=1
M422 427 983 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=144130 $D=1
M423 422 416 425 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=134870 $D=1
M424 423 417 426 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=139500 $D=1
M425 424 418 427 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=144130 $D=1
M426 425 56 242 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=134870 $D=1
M427 426 56 243 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=139500 $D=1
M428 427 56 244 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=144130 $D=1
M429 248 57 425 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=134870 $D=1
M430 249 57 426 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=139500 $D=1
M431 250 57 427 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=144130 $D=1
M432 428 57 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=134870 $D=1
M433 429 57 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=139500 $D=1
M434 430 57 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=144130 $D=1
M435 8 58 431 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=134870 $D=1
M436 9 58 432 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=139500 $D=1
M437 136 58 433 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=144130 $D=1
M438 434 59 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=134870 $D=1
M439 435 59 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=139500 $D=1
M440 436 59 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=144130 $D=1
M441 437 58 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=134870 $D=1
M442 438 58 228 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=139500 $D=1
M443 439 58 229 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=144130 $D=1
M444 8 437 984 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=134870 $D=1
M445 9 438 985 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=139500 $D=1
M446 136 439 986 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=144130 $D=1
M447 440 984 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=134870 $D=1
M448 441 985 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=139500 $D=1
M449 442 986 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=144130 $D=1
M450 437 431 440 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=134870 $D=1
M451 438 432 441 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=139500 $D=1
M452 439 433 442 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=144130 $D=1
M453 440 59 242 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=134870 $D=1
M454 441 59 243 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=139500 $D=1
M455 442 59 244 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=144130 $D=1
M456 248 60 440 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=134870 $D=1
M457 249 60 441 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=139500 $D=1
M458 250 60 442 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=144130 $D=1
M459 443 60 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=134870 $D=1
M460 444 60 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=139500 $D=1
M461 445 60 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=144130 $D=1
M462 8 61 446 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=134870 $D=1
M463 9 61 447 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=139500 $D=1
M464 136 61 448 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=144130 $D=1
M465 449 62 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=134870 $D=1
M466 450 62 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=139500 $D=1
M467 451 62 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=144130 $D=1
M468 452 61 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=134870 $D=1
M469 453 61 228 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=139500 $D=1
M470 454 61 229 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=144130 $D=1
M471 8 452 987 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=134870 $D=1
M472 9 453 988 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=139500 $D=1
M473 136 454 989 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=144130 $D=1
M474 455 987 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=134870 $D=1
M475 456 988 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=139500 $D=1
M476 457 989 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=144130 $D=1
M477 452 446 455 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=134870 $D=1
M478 453 447 456 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=139500 $D=1
M479 454 448 457 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=144130 $D=1
M480 455 62 242 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=134870 $D=1
M481 456 62 243 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=139500 $D=1
M482 457 62 244 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=144130 $D=1
M483 248 63 455 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=134870 $D=1
M484 249 63 456 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=139500 $D=1
M485 250 63 457 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=144130 $D=1
M486 458 63 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=134870 $D=1
M487 459 63 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=139500 $D=1
M488 460 63 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=144130 $D=1
M489 8 64 461 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=134870 $D=1
M490 9 64 462 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=139500 $D=1
M491 136 64 463 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=144130 $D=1
M492 464 65 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=134870 $D=1
M493 465 65 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=139500 $D=1
M494 466 65 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=144130 $D=1
M495 467 64 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=134870 $D=1
M496 468 64 228 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=139500 $D=1
M497 469 64 229 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=144130 $D=1
M498 8 467 990 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=134870 $D=1
M499 9 468 991 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=139500 $D=1
M500 136 469 992 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=144130 $D=1
M501 470 990 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=134870 $D=1
M502 471 991 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=139500 $D=1
M503 472 992 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=144130 $D=1
M504 467 461 470 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=134870 $D=1
M505 468 462 471 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=139500 $D=1
M506 469 463 472 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=144130 $D=1
M507 470 65 242 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=134870 $D=1
M508 471 65 243 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=139500 $D=1
M509 472 65 244 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=144130 $D=1
M510 248 66 470 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=134870 $D=1
M511 249 66 471 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=139500 $D=1
M512 250 66 472 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=144130 $D=1
M513 473 66 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=134870 $D=1
M514 474 66 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=139500 $D=1
M515 475 66 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=144130 $D=1
M516 8 67 476 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=134870 $D=1
M517 9 67 477 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=139500 $D=1
M518 136 67 478 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=144130 $D=1
M519 479 68 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=134870 $D=1
M520 480 68 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=139500 $D=1
M521 481 68 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=144130 $D=1
M522 482 67 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=134870 $D=1
M523 483 67 228 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=139500 $D=1
M524 484 67 229 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=144130 $D=1
M525 8 482 993 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=134870 $D=1
M526 9 483 994 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=139500 $D=1
M527 136 484 995 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=144130 $D=1
M528 485 993 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=134870 $D=1
M529 486 994 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=139500 $D=1
M530 487 995 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=144130 $D=1
M531 482 476 485 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=134870 $D=1
M532 483 477 486 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=139500 $D=1
M533 484 478 487 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=144130 $D=1
M534 485 68 242 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=134870 $D=1
M535 486 68 243 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=139500 $D=1
M536 487 68 244 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=144130 $D=1
M537 248 69 485 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=134870 $D=1
M538 249 69 486 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=139500 $D=1
M539 250 69 487 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=144130 $D=1
M540 488 69 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=134870 $D=1
M541 489 69 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=139500 $D=1
M542 490 69 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=144130 $D=1
M543 8 70 491 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=134870 $D=1
M544 9 70 492 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=139500 $D=1
M545 136 70 493 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=144130 $D=1
M546 494 71 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=134870 $D=1
M547 495 71 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=139500 $D=1
M548 496 71 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=144130 $D=1
M549 497 70 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=134870 $D=1
M550 498 70 228 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=139500 $D=1
M551 499 70 229 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=144130 $D=1
M552 8 497 996 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=134870 $D=1
M553 9 498 997 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=139500 $D=1
M554 136 499 998 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=144130 $D=1
M555 500 996 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=134870 $D=1
M556 501 997 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=139500 $D=1
M557 502 998 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=144130 $D=1
M558 497 491 500 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=134870 $D=1
M559 498 492 501 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=139500 $D=1
M560 499 493 502 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=144130 $D=1
M561 500 71 242 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=134870 $D=1
M562 501 71 243 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=139500 $D=1
M563 502 71 244 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=144130 $D=1
M564 248 72 500 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=134870 $D=1
M565 249 72 501 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=139500 $D=1
M566 250 72 502 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=144130 $D=1
M567 503 72 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=134870 $D=1
M568 504 72 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=139500 $D=1
M569 505 72 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=144130 $D=1
M570 8 73 506 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=134870 $D=1
M571 9 73 507 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=139500 $D=1
M572 136 73 508 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=144130 $D=1
M573 509 74 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=134870 $D=1
M574 510 74 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=139500 $D=1
M575 511 74 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=144130 $D=1
M576 512 73 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=134870 $D=1
M577 513 73 228 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=139500 $D=1
M578 514 73 229 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=144130 $D=1
M579 8 512 999 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=134870 $D=1
M580 9 513 1000 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=139500 $D=1
M581 136 514 1001 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=144130 $D=1
M582 515 999 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=134870 $D=1
M583 516 1000 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=139500 $D=1
M584 517 1001 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=144130 $D=1
M585 512 506 515 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=134870 $D=1
M586 513 507 516 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=139500 $D=1
M587 514 508 517 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=144130 $D=1
M588 515 74 242 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=134870 $D=1
M589 516 74 243 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=139500 $D=1
M590 517 74 244 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=144130 $D=1
M591 248 75 515 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=134870 $D=1
M592 249 75 516 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=139500 $D=1
M593 250 75 517 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=144130 $D=1
M594 518 75 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=134870 $D=1
M595 519 75 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=139500 $D=1
M596 520 75 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=144130 $D=1
M597 8 76 521 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=134870 $D=1
M598 9 76 522 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=139500 $D=1
M599 136 76 523 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=144130 $D=1
M600 524 77 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=134870 $D=1
M601 525 77 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=139500 $D=1
M602 526 77 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=144130 $D=1
M603 527 76 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=134870 $D=1
M604 528 76 228 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=139500 $D=1
M605 529 76 229 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=144130 $D=1
M606 8 527 1002 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=134870 $D=1
M607 9 528 1003 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=139500 $D=1
M608 136 529 1004 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=144130 $D=1
M609 530 1002 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=134870 $D=1
M610 531 1003 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=139500 $D=1
M611 532 1004 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=144130 $D=1
M612 527 521 530 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=134870 $D=1
M613 528 522 531 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=139500 $D=1
M614 529 523 532 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=144130 $D=1
M615 530 77 242 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=134870 $D=1
M616 531 77 243 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=139500 $D=1
M617 532 77 244 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=144130 $D=1
M618 248 78 530 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=134870 $D=1
M619 249 78 531 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=139500 $D=1
M620 250 78 532 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=144130 $D=1
M621 533 78 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=134870 $D=1
M622 534 78 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=139500 $D=1
M623 535 78 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=144130 $D=1
M624 8 79 536 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=134870 $D=1
M625 9 79 537 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=139500 $D=1
M626 136 79 538 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=144130 $D=1
M627 539 80 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=134870 $D=1
M628 540 80 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=139500 $D=1
M629 541 80 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=144130 $D=1
M630 542 79 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=134870 $D=1
M631 543 79 228 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=139500 $D=1
M632 544 79 229 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=144130 $D=1
M633 8 542 1005 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=134870 $D=1
M634 9 543 1006 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=139500 $D=1
M635 136 544 1007 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=144130 $D=1
M636 545 1005 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=134870 $D=1
M637 546 1006 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=139500 $D=1
M638 547 1007 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=144130 $D=1
M639 542 536 545 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=134870 $D=1
M640 543 537 546 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=139500 $D=1
M641 544 538 547 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=144130 $D=1
M642 545 80 242 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=134870 $D=1
M643 546 80 243 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=139500 $D=1
M644 547 80 244 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=144130 $D=1
M645 248 81 545 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=134870 $D=1
M646 249 81 546 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=139500 $D=1
M647 250 81 547 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=144130 $D=1
M648 548 81 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=134870 $D=1
M649 549 81 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=139500 $D=1
M650 550 81 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=144130 $D=1
M651 8 82 551 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=134870 $D=1
M652 9 82 552 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=139500 $D=1
M653 136 82 553 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=144130 $D=1
M654 554 83 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=134870 $D=1
M655 555 83 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=139500 $D=1
M656 556 83 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=144130 $D=1
M657 557 82 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=134870 $D=1
M658 558 82 228 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=139500 $D=1
M659 559 82 229 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=144130 $D=1
M660 8 557 1008 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=134870 $D=1
M661 9 558 1009 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=139500 $D=1
M662 136 559 1010 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=144130 $D=1
M663 560 1008 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=134870 $D=1
M664 561 1009 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=139500 $D=1
M665 562 1010 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=144130 $D=1
M666 557 551 560 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=134870 $D=1
M667 558 552 561 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=139500 $D=1
M668 559 553 562 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=144130 $D=1
M669 560 83 242 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=134870 $D=1
M670 561 83 243 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=139500 $D=1
M671 562 83 244 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=144130 $D=1
M672 248 84 560 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=134870 $D=1
M673 249 84 561 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=139500 $D=1
M674 250 84 562 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=144130 $D=1
M675 563 84 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=134870 $D=1
M676 564 84 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=139500 $D=1
M677 565 84 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=144130 $D=1
M678 8 85 566 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=134870 $D=1
M679 9 85 567 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=139500 $D=1
M680 136 85 568 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=144130 $D=1
M681 569 86 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=134870 $D=1
M682 570 86 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=139500 $D=1
M683 571 86 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=144130 $D=1
M684 572 85 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=134870 $D=1
M685 573 85 228 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=139500 $D=1
M686 574 85 229 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=144130 $D=1
M687 8 572 1011 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=134870 $D=1
M688 9 573 1012 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=139500 $D=1
M689 136 574 1013 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=144130 $D=1
M690 575 1011 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=134870 $D=1
M691 576 1012 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=139500 $D=1
M692 577 1013 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=144130 $D=1
M693 572 566 575 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=134870 $D=1
M694 573 567 576 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=139500 $D=1
M695 574 568 577 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=144130 $D=1
M696 575 86 242 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=134870 $D=1
M697 576 86 243 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=139500 $D=1
M698 577 86 244 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=144130 $D=1
M699 248 87 575 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=134870 $D=1
M700 249 87 576 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=139500 $D=1
M701 250 87 577 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=144130 $D=1
M702 578 87 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=134870 $D=1
M703 579 87 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=139500 $D=1
M704 580 87 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=144130 $D=1
M705 8 88 581 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=134870 $D=1
M706 9 88 582 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=139500 $D=1
M707 136 88 583 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=144130 $D=1
M708 584 89 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=134870 $D=1
M709 585 89 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=139500 $D=1
M710 586 89 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=144130 $D=1
M711 587 88 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=134870 $D=1
M712 588 88 228 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=139500 $D=1
M713 589 88 229 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=144130 $D=1
M714 8 587 1014 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=134870 $D=1
M715 9 588 1015 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=139500 $D=1
M716 136 589 1016 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=144130 $D=1
M717 590 1014 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=134870 $D=1
M718 591 1015 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=139500 $D=1
M719 592 1016 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=144130 $D=1
M720 587 581 590 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=134870 $D=1
M721 588 582 591 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=139500 $D=1
M722 589 583 592 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=144130 $D=1
M723 590 89 242 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=134870 $D=1
M724 591 89 243 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=139500 $D=1
M725 592 89 244 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=144130 $D=1
M726 248 90 590 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=134870 $D=1
M727 249 90 591 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=139500 $D=1
M728 250 90 592 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=144130 $D=1
M729 593 90 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=134870 $D=1
M730 594 90 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=139500 $D=1
M731 595 90 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=144130 $D=1
M732 8 91 596 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=134870 $D=1
M733 9 91 597 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=139500 $D=1
M734 136 91 598 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=144130 $D=1
M735 599 92 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=134870 $D=1
M736 600 92 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=139500 $D=1
M737 601 92 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=144130 $D=1
M738 602 91 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=134870 $D=1
M739 603 91 228 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=139500 $D=1
M740 604 91 229 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=144130 $D=1
M741 8 602 1017 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=134870 $D=1
M742 9 603 1018 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=139500 $D=1
M743 136 604 1019 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=144130 $D=1
M744 605 1017 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=134870 $D=1
M745 606 1018 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=139500 $D=1
M746 607 1019 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=144130 $D=1
M747 602 596 605 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=134870 $D=1
M748 603 597 606 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=139500 $D=1
M749 604 598 607 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=144130 $D=1
M750 605 92 242 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=134870 $D=1
M751 606 92 243 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=139500 $D=1
M752 607 92 244 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=144130 $D=1
M753 248 93 605 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=134870 $D=1
M754 249 93 606 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=139500 $D=1
M755 250 93 607 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=144130 $D=1
M756 608 93 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=134870 $D=1
M757 609 93 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=139500 $D=1
M758 610 93 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=144130 $D=1
M759 8 94 611 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=134870 $D=1
M760 9 94 612 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=139500 $D=1
M761 136 94 613 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=144130 $D=1
M762 614 95 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=134870 $D=1
M763 615 95 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=139500 $D=1
M764 616 95 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=144130 $D=1
M765 617 94 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=134870 $D=1
M766 618 94 228 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=139500 $D=1
M767 619 94 229 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=144130 $D=1
M768 8 617 1020 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=134870 $D=1
M769 9 618 1021 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=139500 $D=1
M770 136 619 1022 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=144130 $D=1
M771 620 1020 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=134870 $D=1
M772 621 1021 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=139500 $D=1
M773 622 1022 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=144130 $D=1
M774 617 611 620 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=134870 $D=1
M775 618 612 621 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=139500 $D=1
M776 619 613 622 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=144130 $D=1
M777 620 95 242 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=134870 $D=1
M778 621 95 243 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=139500 $D=1
M779 622 95 244 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=144130 $D=1
M780 248 96 620 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=134870 $D=1
M781 249 96 621 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=139500 $D=1
M782 250 96 622 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=144130 $D=1
M783 623 96 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=134870 $D=1
M784 624 96 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=139500 $D=1
M785 625 96 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=144130 $D=1
M786 8 97 626 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=134870 $D=1
M787 9 97 627 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=139500 $D=1
M788 136 97 628 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=144130 $D=1
M789 629 98 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=134870 $D=1
M790 630 98 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=139500 $D=1
M791 631 98 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=144130 $D=1
M792 632 97 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=134870 $D=1
M793 633 97 228 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=139500 $D=1
M794 634 97 229 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=144130 $D=1
M795 8 632 1023 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=134870 $D=1
M796 9 633 1024 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=139500 $D=1
M797 136 634 1025 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=144130 $D=1
M798 635 1023 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=134870 $D=1
M799 636 1024 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=139500 $D=1
M800 637 1025 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=144130 $D=1
M801 632 626 635 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=134870 $D=1
M802 633 627 636 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=139500 $D=1
M803 634 628 637 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=144130 $D=1
M804 635 98 242 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=134870 $D=1
M805 636 98 243 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=139500 $D=1
M806 637 98 244 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=144130 $D=1
M807 248 99 635 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=134870 $D=1
M808 249 99 636 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=139500 $D=1
M809 250 99 637 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=144130 $D=1
M810 638 99 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=134870 $D=1
M811 639 99 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=139500 $D=1
M812 640 99 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=144130 $D=1
M813 8 100 641 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=134870 $D=1
M814 9 100 642 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=139500 $D=1
M815 136 100 643 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=144130 $D=1
M816 644 101 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=134870 $D=1
M817 645 101 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=139500 $D=1
M818 646 101 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=144130 $D=1
M819 647 100 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=134870 $D=1
M820 648 100 228 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=139500 $D=1
M821 649 100 229 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=144130 $D=1
M822 8 647 1026 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=134870 $D=1
M823 9 648 1027 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=139500 $D=1
M824 136 649 1028 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=144130 $D=1
M825 650 1026 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=134870 $D=1
M826 651 1027 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=139500 $D=1
M827 652 1028 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=144130 $D=1
M828 647 641 650 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=134870 $D=1
M829 648 642 651 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=139500 $D=1
M830 649 643 652 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=144130 $D=1
M831 650 101 242 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=134870 $D=1
M832 651 101 243 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=139500 $D=1
M833 652 101 244 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=144130 $D=1
M834 248 102 650 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=134870 $D=1
M835 249 102 651 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=139500 $D=1
M836 250 102 652 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=144130 $D=1
M837 653 102 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=134870 $D=1
M838 654 102 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=139500 $D=1
M839 655 102 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=144130 $D=1
M840 8 103 656 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=134870 $D=1
M841 9 103 657 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=139500 $D=1
M842 136 103 658 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=144130 $D=1
M843 659 104 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=134870 $D=1
M844 660 104 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=139500 $D=1
M845 661 104 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=144130 $D=1
M846 662 103 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=134870 $D=1
M847 663 103 228 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=139500 $D=1
M848 664 103 229 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=144130 $D=1
M849 8 662 1029 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=134870 $D=1
M850 9 663 1030 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=139500 $D=1
M851 136 664 1031 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=144130 $D=1
M852 665 1029 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=134870 $D=1
M853 666 1030 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=139500 $D=1
M854 667 1031 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=144130 $D=1
M855 662 656 665 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=134870 $D=1
M856 663 657 666 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=139500 $D=1
M857 664 658 667 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=144130 $D=1
M858 665 104 242 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=134870 $D=1
M859 666 104 243 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=139500 $D=1
M860 667 104 244 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=144130 $D=1
M861 248 105 665 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=134870 $D=1
M862 249 105 666 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=139500 $D=1
M863 250 105 667 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=144130 $D=1
M864 668 105 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=134870 $D=1
M865 669 105 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=139500 $D=1
M866 670 105 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=144130 $D=1
M867 8 106 671 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=134870 $D=1
M868 9 106 672 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=139500 $D=1
M869 136 106 673 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=144130 $D=1
M870 674 107 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=134870 $D=1
M871 675 107 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=139500 $D=1
M872 676 107 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=144130 $D=1
M873 677 106 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=134870 $D=1
M874 678 106 228 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=139500 $D=1
M875 679 106 229 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=144130 $D=1
M876 8 677 1032 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=134870 $D=1
M877 9 678 1033 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=139500 $D=1
M878 136 679 1034 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=144130 $D=1
M879 680 1032 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=134870 $D=1
M880 681 1033 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=139500 $D=1
M881 682 1034 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=144130 $D=1
M882 677 671 680 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=134870 $D=1
M883 678 672 681 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=139500 $D=1
M884 679 673 682 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=144130 $D=1
M885 680 107 242 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=134870 $D=1
M886 681 107 243 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=139500 $D=1
M887 682 107 244 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=144130 $D=1
M888 248 108 680 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=134870 $D=1
M889 249 108 681 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=139500 $D=1
M890 250 108 682 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=144130 $D=1
M891 683 108 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=134870 $D=1
M892 684 108 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=139500 $D=1
M893 685 108 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=144130 $D=1
M894 8 109 686 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=134870 $D=1
M895 9 109 687 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=139500 $D=1
M896 136 109 688 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=144130 $D=1
M897 689 110 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=134870 $D=1
M898 690 110 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=139500 $D=1
M899 691 110 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=144130 $D=1
M900 692 109 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=134870 $D=1
M901 693 109 228 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=139500 $D=1
M902 694 109 229 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=144130 $D=1
M903 8 692 1035 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=134870 $D=1
M904 9 693 1036 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=139500 $D=1
M905 136 694 1037 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=144130 $D=1
M906 695 1035 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=134870 $D=1
M907 696 1036 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=139500 $D=1
M908 697 1037 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=144130 $D=1
M909 692 686 695 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=134870 $D=1
M910 693 687 696 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=139500 $D=1
M911 694 688 697 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=144130 $D=1
M912 695 110 242 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=134870 $D=1
M913 696 110 243 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=139500 $D=1
M914 697 110 244 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=144130 $D=1
M915 248 111 695 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=134870 $D=1
M916 249 111 696 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=139500 $D=1
M917 250 111 697 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=144130 $D=1
M918 698 111 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=134870 $D=1
M919 699 111 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=139500 $D=1
M920 700 111 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=144130 $D=1
M921 8 112 701 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=134870 $D=1
M922 9 112 702 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=139500 $D=1
M923 136 112 703 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=144130 $D=1
M924 704 113 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=134870 $D=1
M925 705 113 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=139500 $D=1
M926 706 113 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=144130 $D=1
M927 8 113 242 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=134870 $D=1
M928 9 113 243 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=139500 $D=1
M929 136 113 244 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=144130 $D=1
M930 248 112 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=134870 $D=1
M931 249 112 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=139500 $D=1
M932 250 112 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=144130 $D=1
M933 8 710 707 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=134870 $D=1
M934 9 711 708 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=139500 $D=1
M935 136 712 709 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=144130 $D=1
M936 710 114 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=134870 $D=1
M937 711 114 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=139500 $D=1
M938 712 114 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=144130 $D=1
M939 1038 242 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=134870 $D=1
M940 1039 243 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=139500 $D=1
M941 1040 244 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=144130 $D=1
M942 713 707 1038 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=134870 $D=1
M943 714 708 1039 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=139500 $D=1
M944 715 709 1040 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=144130 $D=1
M945 8 713 716 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=134870 $D=1
M946 9 714 717 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=139500 $D=1
M947 136 715 718 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=144130 $D=1
M948 1041 716 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=134870 $D=1
M949 1042 717 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=139500 $D=1
M950 1043 718 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=144130 $D=1
M951 713 710 1041 8 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=134870 $D=1
M952 714 711 1042 9 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=139500 $D=1
M953 715 712 1043 136 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=144130 $D=1
M954 8 722 719 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=134870 $D=1
M955 9 723 720 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=139500 $D=1
M956 136 724 721 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=144130 $D=1
M957 722 114 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=134870 $D=1
M958 723 114 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=139500 $D=1
M959 724 114 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=144130 $D=1
M960 1044 248 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=134870 $D=1
M961 1045 249 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=139500 $D=1
M962 1046 250 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=144130 $D=1
M963 725 719 1044 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=134870 $D=1
M964 726 720 1045 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=139500 $D=1
M965 727 721 1046 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=144130 $D=1
M966 8 725 115 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=134870 $D=1
M967 9 726 116 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=139500 $D=1
M968 136 727 117 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=144130 $D=1
M969 1047 115 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=134870 $D=1
M970 1048 116 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=139500 $D=1
M971 1049 117 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=144130 $D=1
M972 725 722 1047 8 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=134870 $D=1
M973 726 723 1048 9 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=139500 $D=1
M974 727 724 1049 136 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=144130 $D=1
M975 728 118 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=134870 $D=1
M976 729 118 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=139500 $D=1
M977 730 118 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=144130 $D=1
M978 731 728 716 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=134870 $D=1
M979 732 729 717 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=139500 $D=1
M980 733 730 718 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=144130 $D=1
M981 119 118 731 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=134870 $D=1
M982 120 118 732 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=139500 $D=1
M983 121 118 733 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=144130 $D=1
M984 734 122 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=134870 $D=1
M985 735 122 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=139500 $D=1
M986 736 122 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=144130 $D=1
M987 737 734 115 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=134870 $D=1
M988 738 735 116 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=139500 $D=1
M989 739 736 117 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=144130 $D=1
M990 1050 122 737 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=134870 $D=1
M991 1051 122 738 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=139500 $D=1
M992 1052 122 739 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=144130 $D=1
M993 8 115 1050 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=134870 $D=1
M994 9 116 1051 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=139500 $D=1
M995 136 117 1052 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=144130 $D=1
M996 740 123 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=134870 $D=1
M997 741 123 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=139500 $D=1
M998 742 123 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=144130 $D=1
M999 124 740 737 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=134870 $D=1
M1000 125 741 738 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=139500 $D=1
M1001 126 742 739 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=144130 $D=1
M1002 11 123 124 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=134870 $D=1
M1003 12 123 125 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=139500 $D=1
M1004 13 123 126 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=144130 $D=1
M1005 745 743 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=134870 $D=1
M1006 746 744 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=139500 $D=1
M1007 747 127 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=144130 $D=1
M1008 8 751 748 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=134870 $D=1
M1009 9 752 749 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=139500 $D=1
M1010 136 753 750 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=144130 $D=1
M1011 754 731 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=134870 $D=1
M1012 755 732 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=139500 $D=1
M1013 756 733 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=144130 $D=1
M1014 751 754 743 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=134870 $D=1
M1015 752 755 744 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=139500 $D=1
M1016 753 756 127 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=144130 $D=1
M1017 745 731 751 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=134870 $D=1
M1018 746 732 752 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=139500 $D=1
M1019 747 733 753 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=144130 $D=1
M1020 757 748 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=134870 $D=1
M1021 758 749 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=139500 $D=1
M1022 759 750 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=144130 $D=1
M1023 128 757 124 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=134870 $D=1
M1024 743 758 125 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=139500 $D=1
M1025 744 759 126 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=144130 $D=1
M1026 731 748 128 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=134870 $D=1
M1027 732 749 743 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=139500 $D=1
M1028 733 750 744 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=144130 $D=1
M1029 760 128 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=134870 $D=1
M1030 761 743 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=139500 $D=1
M1031 762 744 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=144130 $D=1
M1032 763 748 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=134870 $D=1
M1033 764 749 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=139500 $D=1
M1034 765 750 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=144130 $D=1
M1035 766 763 760 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=134870 $D=1
M1036 767 764 761 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=139500 $D=1
M1037 768 765 762 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=144130 $D=1
M1038 124 748 766 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=134870 $D=1
M1039 125 749 767 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=139500 $D=1
M1040 126 750 768 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=144130 $D=1
M1041 769 731 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=134870 $D=1
M1042 770 732 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=139500 $D=1
M1043 771 733 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=144130 $D=1
M1044 8 124 769 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=134870 $D=1
M1045 9 125 770 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=139500 $D=1
M1046 136 126 771 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=144130 $D=1
M1047 772 766 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=134870 $D=1
M1048 773 767 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=139500 $D=1
M1049 774 768 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=144130 $D=1
M1050 1092 731 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=134870 $D=1
M1051 1093 732 9 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=139500 $D=1
M1052 1094 733 136 136 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=144130 $D=1
M1053 775 124 1092 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=134870 $D=1
M1054 776 125 1093 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=139500 $D=1
M1055 777 126 1094 136 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=144130 $D=1
M1056 1095 731 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=134870 $D=1
M1057 1096 732 9 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=139500 $D=1
M1058 1097 733 136 136 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=144130 $D=1
M1059 778 124 1095 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=134870 $D=1
M1060 779 125 1096 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=139500 $D=1
M1061 780 126 1097 136 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=144130 $D=1
M1062 784 731 781 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=134870 $D=1
M1063 785 732 782 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=139500 $D=1
M1064 786 733 783 136 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=144130 $D=1
M1065 781 124 784 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=134870 $D=1
M1066 782 125 785 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=139500 $D=1
M1067 783 126 786 136 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=144130 $D=1
M1068 8 778 781 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=134870 $D=1
M1069 9 779 782 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=139500 $D=1
M1070 136 780 783 136 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=144130 $D=1
M1071 787 132 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=134870 $D=1
M1072 788 132 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=139500 $D=1
M1073 789 132 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=144130 $D=1
M1074 790 787 769 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=134870 $D=1
M1075 791 788 770 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=139500 $D=1
M1076 792 789 771 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=144130 $D=1
M1077 775 132 790 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=134870 $D=1
M1078 776 132 791 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=139500 $D=1
M1079 777 132 792 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=144130 $D=1
M1080 793 787 772 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=134870 $D=1
M1081 794 788 773 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=139500 $D=1
M1082 795 789 774 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=144130 $D=1
M1083 784 132 793 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=134870 $D=1
M1084 785 132 794 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=139500 $D=1
M1085 786 132 795 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=144130 $D=1
M1086 796 133 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=134870 $D=1
M1087 797 133 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=139500 $D=1
M1088 798 133 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=144130 $D=1
M1089 799 796 793 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=134870 $D=1
M1090 800 797 794 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=139500 $D=1
M1091 801 798 795 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=144130 $D=1
M1092 790 133 799 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=134870 $D=1
M1093 791 133 800 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=139500 $D=1
M1094 792 133 801 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=144130 $D=1
M1095 14 799 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=134870 $D=1
M1096 15 800 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=139500 $D=1
M1097 16 801 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=144130 $D=1
M1098 802 134 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=134870 $D=1
M1099 803 134 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=139500 $D=1
M1100 804 134 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=144130 $D=1
M1101 805 802 125 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=134870 $D=1
M1102 806 803 135 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=139500 $D=1
M1103 807 804 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=144130 $D=1
M1104 137 134 805 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=134870 $D=1
M1105 124 134 806 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=139500 $D=1
M1106 125 134 807 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=144130 $D=1
M1107 808 134 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=134870 $D=1
M1108 809 134 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=139500 $D=1
M1109 810 134 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=144130 $D=1
M1110 817 808 138 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=134870 $D=1
M1111 818 809 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=139500 $D=1
M1112 819 810 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=144130 $D=1
M1113 139 134 817 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=134870 $D=1
M1114 140 134 818 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=139500 $D=1
M1115 141 134 819 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=144130 $D=1
M1116 820 134 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=134870 $D=1
M1117 821 134 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=139500 $D=1
M1118 822 134 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=144130 $D=1
M1119 823 820 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=134870 $D=1
M1120 824 821 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=139500 $D=1
M1121 825 822 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=144130 $D=1
M1122 142 134 823 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=134870 $D=1
M1123 143 134 824 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=139500 $D=1
M1124 144 134 825 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=144130 $D=1
M1125 826 134 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=134870 $D=1
M1126 827 134 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=139500 $D=1
M1127 828 134 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=144130 $D=1
M1128 829 826 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=134870 $D=1
M1129 830 827 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=139500 $D=1
M1130 831 828 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=144130 $D=1
M1131 145 134 829 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=134870 $D=1
M1132 146 134 830 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=139500 $D=1
M1133 147 134 831 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=144130 $D=1
M1134 832 134 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=134870 $D=1
M1135 833 134 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=139500 $D=1
M1136 834 134 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=144130 $D=1
M1137 835 832 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=134870 $D=1
M1138 836 833 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=139500 $D=1
M1139 837 834 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=144130 $D=1
M1140 148 134 835 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=134870 $D=1
M1141 149 134 836 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=139500 $D=1
M1142 144 134 837 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=144130 $D=1
M1143 8 731 1065 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=134870 $D=1
M1144 9 732 1066 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=139500 $D=1
M1145 136 733 1067 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=144130 $D=1
M1146 124 1065 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=134870 $D=1
M1147 125 1066 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=139500 $D=1
M1148 135 1067 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=144130 $D=1
M1149 838 126 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=134870 $D=1
M1150 839 126 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=139500 $D=1
M1151 840 126 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=144130 $D=1
M1152 141 838 124 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=134870 $D=1
M1153 150 839 125 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=139500 $D=1
M1154 138 840 135 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=144130 $D=1
M1155 805 126 141 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=134870 $D=1
M1156 806 126 150 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=139500 $D=1
M1157 807 126 138 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=144130 $D=1
M1158 841 125 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=134870 $D=1
M1159 842 125 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=139500 $D=1
M1160 843 125 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=144130 $D=1
M1161 131 841 141 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=134870 $D=1
M1162 130 842 150 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=139500 $D=1
M1163 129 843 138 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=144130 $D=1
M1164 817 125 131 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=134870 $D=1
M1165 818 125 130 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=139500 $D=1
M1166 819 125 129 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=144130 $D=1
M1167 844 124 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=134870 $D=1
M1168 845 124 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=139500 $D=1
M1169 846 124 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=144130 $D=1
M1170 151 844 131 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=134870 $D=1
M1171 152 845 130 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=139500 $D=1
M1172 153 846 129 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=144130 $D=1
M1173 823 124 151 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=134870 $D=1
M1174 824 124 152 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=139500 $D=1
M1175 825 124 153 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=144130 $D=1
M1176 847 154 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=134870 $D=1
M1177 848 154 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=139500 $D=1
M1178 849 154 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=144130 $D=1
M1179 155 847 151 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=134870 $D=1
M1180 156 848 152 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=139500 $D=1
M1181 157 849 153 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=144130 $D=1
M1182 829 154 155 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=134870 $D=1
M1183 830 154 156 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=139500 $D=1
M1184 831 154 157 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=144130 $D=1
M1185 850 158 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=134870 $D=1
M1186 851 158 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=139500 $D=1
M1187 852 158 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=144130 $D=1
M1188 206 850 155 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=134870 $D=1
M1189 207 851 156 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=139500 $D=1
M1190 208 852 157 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=144130 $D=1
M1191 835 158 206 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=134870 $D=1
M1192 836 158 207 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=139500 $D=1
M1193 837 158 208 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=144130 $D=1
M1194 853 159 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=134870 $D=1
M1195 854 159 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=139500 $D=1
M1196 855 159 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=144130 $D=1
M1197 856 853 115 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=134870 $D=1
M1198 857 854 116 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=139500 $D=1
M1199 858 855 117 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=144130 $D=1
M1200 11 159 856 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=134870 $D=1
M1201 12 159 857 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=139500 $D=1
M1202 13 159 858 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=144130 $D=1
M1203 1098 716 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=134870 $D=1
M1204 1099 717 9 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=139500 $D=1
M1205 1100 718 136 136 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=144130 $D=1
M1206 859 856 1098 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=134870 $D=1
M1207 860 857 1099 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=139500 $D=1
M1208 861 858 1100 136 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=144130 $D=1
M1209 865 716 862 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=134870 $D=1
M1210 866 717 863 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=139500 $D=1
M1211 867 718 864 136 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=144130 $D=1
M1212 862 856 865 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=134870 $D=1
M1213 863 857 866 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=139500 $D=1
M1214 864 858 867 136 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=144130 $D=1
M1215 8 859 862 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=134870 $D=1
M1216 9 860 863 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=139500 $D=1
M1217 136 861 864 136 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=144130 $D=1
M1218 1101 868 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=134870 $D=1
M1219 1102 869 9 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=139500 $D=1
M1220 1103 870 136 136 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=144130 $D=1
M1221 1068 865 1101 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=134870 $D=1
M1222 1069 866 1102 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=139500 $D=1
M1223 1070 867 1103 136 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=144130 $D=1
M1224 869 1068 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=134870 $D=1
M1225 871 1069 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=139500 $D=1
M1226 160 1070 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=144130 $D=1
M1227 872 716 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=134870 $D=1
M1228 873 717 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=139500 $D=1
M1229 874 718 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=144130 $D=1
M1230 8 875 872 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=134870 $D=1
M1231 9 876 873 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=139500 $D=1
M1232 136 877 874 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=144130 $D=1
M1233 875 856 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=134870 $D=1
M1234 876 857 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=139500 $D=1
M1235 877 858 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=144130 $D=1
M1236 1104 872 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=134870 $D=1
M1237 1105 873 9 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=139500 $D=1
M1238 1106 874 136 136 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=144130 $D=1
M1239 878 868 1104 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=134870 $D=1
M1240 879 869 1105 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=139500 $D=1
M1241 880 870 1106 136 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=144130 $D=1
M1242 883 161 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=134870 $D=1
M1243 884 881 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=139500 $D=1
M1244 885 882 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=144130 $D=1
M1245 1107 878 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=134870 $D=1
M1246 1108 879 9 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=139500 $D=1
M1247 1109 880 136 136 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=144130 $D=1
M1248 881 883 1107 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=134870 $D=1
M1249 882 884 1108 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=139500 $D=1
M1250 162 885 1109 136 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=144130 $D=1
M1251 888 886 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=134870 $D=1
M1252 889 887 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=139500 $D=1
M1253 890 136 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=144130 $D=1
M1254 8 894 891 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=134870 $D=1
M1255 9 895 892 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=139500 $D=1
M1256 136 896 893 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=144130 $D=1
M1257 897 119 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=134870 $D=1
M1258 898 120 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=139500 $D=1
M1259 899 121 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=144130 $D=1
M1260 894 897 886 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=134870 $D=1
M1261 895 898 887 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=139500 $D=1
M1262 896 899 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=144130 $D=1
M1263 888 119 894 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=134870 $D=1
M1264 889 120 895 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=139500 $D=1
M1265 890 121 896 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=144130 $D=1
M1266 900 891 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=134870 $D=1
M1267 901 892 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=139500 $D=1
M1268 902 893 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=144130 $D=1
M1269 164 900 163 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=134870 $D=1
M1270 886 901 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=139500 $D=1
M1271 887 902 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=144130 $D=1
M1272 119 891 164 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=134870 $D=1
M1273 120 892 886 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=139500 $D=1
M1274 121 893 887 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=144130 $D=1
M1275 903 164 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=134870 $D=1
M1276 904 886 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=139500 $D=1
M1277 905 887 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=144130 $D=1
M1278 906 891 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=134870 $D=1
M1279 907 892 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=139500 $D=1
M1280 908 893 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=144130 $D=1
M1281 209 906 903 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=134870 $D=1
M1282 210 907 904 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=139500 $D=1
M1283 211 908 905 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=144130 $D=1
M1284 163 891 209 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=134870 $D=1
M1285 9 892 210 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=139500 $D=1
M1286 136 893 211 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=144130 $D=1
M1287 909 165 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=134870 $D=1
M1288 910 165 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=139500 $D=1
M1289 911 165 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=144130 $D=1
M1290 912 909 209 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=134870 $D=1
M1291 913 910 210 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=139500 $D=1
M1292 914 911 211 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=144130 $D=1
M1293 14 165 912 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=134870 $D=1
M1294 15 165 913 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=139500 $D=1
M1295 16 165 914 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=144130 $D=1
M1296 915 166 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=134870 $D=1
M1297 916 166 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=139500 $D=1
M1298 917 166 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=144130 $D=1
M1299 166 915 912 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=134870 $D=1
M1300 166 916 913 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=139500 $D=1
M1301 166 917 914 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=144130 $D=1
M1302 8 166 166 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=134870 $D=1
M1303 9 166 166 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=139500 $D=1
M1304 136 166 166 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=144130 $D=1
M1305 918 114 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=134870 $D=1
M1306 919 114 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=139500 $D=1
M1307 920 114 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=144130 $D=1
M1308 8 918 921 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=134870 $D=1
M1309 9 919 922 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=139500 $D=1
M1310 136 920 923 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=144130 $D=1
M1311 924 114 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=134870 $D=1
M1312 925 114 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=139500 $D=1
M1313 926 114 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=144130 $D=1
M1314 927 918 166 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=134870 $D=1
M1315 928 919 166 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=139500 $D=1
M1316 929 920 166 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=144130 $D=1
M1317 8 927 1071 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=134870 $D=1
M1318 9 928 1072 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=139500 $D=1
M1319 136 929 1073 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=144130 $D=1
M1320 930 1071 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=134870 $D=1
M1321 931 1072 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=139500 $D=1
M1322 932 1073 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=144130 $D=1
M1323 927 921 930 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=134870 $D=1
M1324 928 922 931 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=139500 $D=1
M1325 929 923 932 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=144130 $D=1
M1326 933 114 930 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=134870 $D=1
M1327 934 114 931 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=139500 $D=1
M1328 935 114 932 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=144130 $D=1
M1329 8 939 936 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=134870 $D=1
M1330 9 940 937 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=139500 $D=1
M1331 136 941 938 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=144130 $D=1
M1332 939 114 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=134870 $D=1
M1333 940 114 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=139500 $D=1
M1334 941 114 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=144130 $D=1
M1335 1074 933 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=134870 $D=1
M1336 1075 934 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=139500 $D=1
M1337 1076 935 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=144130 $D=1
M1338 942 936 1074 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=134870 $D=1
M1339 943 937 1075 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=139500 $D=1
M1340 944 938 1076 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=144130 $D=1
M1341 8 942 119 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=134870 $D=1
M1342 9 943 120 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=139500 $D=1
M1343 136 944 121 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=144130 $D=1
M1344 1077 119 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=134870 $D=1
M1345 1078 120 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=139500 $D=1
M1346 1079 121 136 136 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=144130 $D=1
M1347 942 939 1077 8 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=134870 $D=1
M1348 943 940 1078 9 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=139500 $D=1
M1349 944 941 1079 136 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=144130 $D=1
M1350 170 1 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=136120 $D=0
M1351 171 1 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=140750 $D=0
M1352 172 1 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=145380 $D=0
M1353 173 1 2 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=136120 $D=0
M1354 174 1 3 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=140750 $D=0
M1355 175 1 4 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=145380 $D=0
M1356 8 170 173 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=136120 $D=0
M1357 9 171 174 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=140750 $D=0
M1358 136 172 175 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=145380 $D=0
M1359 176 1 2 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=136120 $D=0
M1360 177 1 3 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=140750 $D=0
M1361 178 1 4 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=145380 $D=0
M1362 2 170 176 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=136120 $D=0
M1363 3 171 177 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=140750 $D=0
M1364 4 172 178 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=145380 $D=0
M1365 179 1 2 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=136120 $D=0
M1366 180 1 3 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=140750 $D=0
M1367 181 1 4 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=145380 $D=0
M1368 2 170 179 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=136120 $D=0
M1369 3 171 180 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=140750 $D=0
M1370 4 172 181 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=145380 $D=0
M1371 185 5 179 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=136120 $D=0
M1372 186 5 180 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=140750 $D=0
M1373 187 5 181 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=145380 $D=0
M1374 182 5 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=136120 $D=0
M1375 183 5 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=140750 $D=0
M1376 184 5 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=145380 $D=0
M1377 188 5 176 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=136120 $D=0
M1378 189 5 177 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=140750 $D=0
M1379 190 5 178 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=145380 $D=0
M1380 173 182 188 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=136120 $D=0
M1381 174 183 189 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=140750 $D=0
M1382 175 184 190 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=145380 $D=0
M1383 191 6 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=136120 $D=0
M1384 192 6 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=140750 $D=0
M1385 193 6 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=145380 $D=0
M1386 194 6 188 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=136120 $D=0
M1387 195 6 189 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=140750 $D=0
M1388 196 6 190 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=145380 $D=0
M1389 185 191 194 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=136120 $D=0
M1390 186 192 195 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=140750 $D=0
M1391 187 193 196 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=145380 $D=0
M1392 197 7 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=136120 $D=0
M1393 198 7 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=140750 $D=0
M1394 199 7 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=145380 $D=0
M1395 200 7 8 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=136120 $D=0
M1396 201 7 9 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=140750 $D=0
M1397 202 7 10 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=145380 $D=0
M1398 11 197 200 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=136120 $D=0
M1399 12 198 201 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=140750 $D=0
M1400 13 199 202 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=145380 $D=0
M1401 203 7 14 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=136120 $D=0
M1402 204 7 15 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=140750 $D=0
M1403 205 7 16 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=145380 $D=0
M1404 206 197 203 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=136120 $D=0
M1405 207 198 204 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=140750 $D=0
M1406 208 199 205 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=145380 $D=0
M1407 212 7 209 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=136120 $D=0
M1408 213 7 210 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=140750 $D=0
M1409 214 7 211 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=145380 $D=0
M1410 194 197 212 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=136120 $D=0
M1411 195 198 213 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=140750 $D=0
M1412 196 199 214 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=145380 $D=0
M1413 218 17 212 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=136120 $D=0
M1414 219 17 213 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=140750 $D=0
M1415 220 17 214 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=145380 $D=0
M1416 215 17 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=136120 $D=0
M1417 216 17 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=140750 $D=0
M1418 217 17 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=145380 $D=0
M1419 221 17 203 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=136120 $D=0
M1420 222 17 204 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=140750 $D=0
M1421 223 17 205 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=145380 $D=0
M1422 200 215 221 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=136120 $D=0
M1423 201 216 222 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=140750 $D=0
M1424 202 217 223 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=145380 $D=0
M1425 224 18 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=136120 $D=0
M1426 225 18 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=140750 $D=0
M1427 226 18 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=145380 $D=0
M1428 227 18 221 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=136120 $D=0
M1429 228 18 222 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=140750 $D=0
M1430 229 18 223 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=145380 $D=0
M1431 218 224 227 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=136120 $D=0
M1432 219 225 228 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=140750 $D=0
M1433 220 226 229 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=145380 $D=0
M1434 163 19 230 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=136120 $D=0
M1435 167 19 231 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=140750 $D=0
M1436 168 19 232 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=145380 $D=0
M1437 233 20 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=136120 $D=0
M1438 234 20 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=140750 $D=0
M1439 235 20 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=145380 $D=0
M1440 236 230 227 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=136120 $D=0
M1441 237 231 228 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=140750 $D=0
M1442 238 232 229 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=145380 $D=0
M1443 163 236 945 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=136120 $D=0
M1444 167 237 946 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=140750 $D=0
M1445 168 238 947 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=145380 $D=0
M1446 239 945 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=136120 $D=0
M1447 240 946 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=140750 $D=0
M1448 241 947 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=145380 $D=0
M1449 236 19 239 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=136120 $D=0
M1450 237 19 240 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=140750 $D=0
M1451 238 19 241 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=145380 $D=0
M1452 239 233 242 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=136120 $D=0
M1453 240 234 243 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=140750 $D=0
M1454 241 235 244 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=145380 $D=0
M1455 248 245 239 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=136120 $D=0
M1456 249 246 240 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=140750 $D=0
M1457 250 247 241 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=145380 $D=0
M1458 245 21 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=136120 $D=0
M1459 246 21 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=140750 $D=0
M1460 247 21 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=145380 $D=0
M1461 163 22 251 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=136120 $D=0
M1462 167 22 252 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=140750 $D=0
M1463 168 22 253 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=145380 $D=0
M1464 254 23 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=136120 $D=0
M1465 255 23 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=140750 $D=0
M1466 256 23 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=145380 $D=0
M1467 257 251 227 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=136120 $D=0
M1468 258 252 228 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=140750 $D=0
M1469 259 253 229 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=145380 $D=0
M1470 163 257 948 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=136120 $D=0
M1471 167 258 949 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=140750 $D=0
M1472 168 259 950 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=145380 $D=0
M1473 260 948 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=136120 $D=0
M1474 261 949 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=140750 $D=0
M1475 262 950 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=145380 $D=0
M1476 257 22 260 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=136120 $D=0
M1477 258 22 261 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=140750 $D=0
M1478 259 22 262 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=145380 $D=0
M1479 260 254 242 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=136120 $D=0
M1480 261 255 243 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=140750 $D=0
M1481 262 256 244 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=145380 $D=0
M1482 248 263 260 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=136120 $D=0
M1483 249 264 261 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=140750 $D=0
M1484 250 265 262 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=145380 $D=0
M1485 263 24 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=136120 $D=0
M1486 264 24 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=140750 $D=0
M1487 265 24 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=145380 $D=0
M1488 163 25 266 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=136120 $D=0
M1489 167 25 267 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=140750 $D=0
M1490 168 25 268 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=145380 $D=0
M1491 269 26 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=136120 $D=0
M1492 270 26 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=140750 $D=0
M1493 271 26 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=145380 $D=0
M1494 272 266 227 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=136120 $D=0
M1495 273 267 228 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=140750 $D=0
M1496 274 268 229 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=145380 $D=0
M1497 163 272 951 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=136120 $D=0
M1498 167 273 952 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=140750 $D=0
M1499 168 274 953 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=145380 $D=0
M1500 275 951 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=136120 $D=0
M1501 276 952 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=140750 $D=0
M1502 277 953 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=145380 $D=0
M1503 272 25 275 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=136120 $D=0
M1504 273 25 276 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=140750 $D=0
M1505 274 25 277 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=145380 $D=0
M1506 275 269 242 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=136120 $D=0
M1507 276 270 243 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=140750 $D=0
M1508 277 271 244 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=145380 $D=0
M1509 248 278 275 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=136120 $D=0
M1510 249 279 276 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=140750 $D=0
M1511 250 280 277 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=145380 $D=0
M1512 278 27 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=136120 $D=0
M1513 279 27 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=140750 $D=0
M1514 280 27 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=145380 $D=0
M1515 163 28 281 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=136120 $D=0
M1516 167 28 282 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=140750 $D=0
M1517 168 28 283 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=145380 $D=0
M1518 284 29 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=136120 $D=0
M1519 285 29 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=140750 $D=0
M1520 286 29 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=145380 $D=0
M1521 287 281 227 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=136120 $D=0
M1522 288 282 228 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=140750 $D=0
M1523 289 283 229 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=145380 $D=0
M1524 163 287 954 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=136120 $D=0
M1525 167 288 955 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=140750 $D=0
M1526 168 289 956 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=145380 $D=0
M1527 290 954 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=136120 $D=0
M1528 291 955 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=140750 $D=0
M1529 292 956 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=145380 $D=0
M1530 287 28 290 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=136120 $D=0
M1531 288 28 291 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=140750 $D=0
M1532 289 28 292 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=145380 $D=0
M1533 290 284 242 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=136120 $D=0
M1534 291 285 243 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=140750 $D=0
M1535 292 286 244 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=145380 $D=0
M1536 248 293 290 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=136120 $D=0
M1537 249 294 291 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=140750 $D=0
M1538 250 295 292 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=145380 $D=0
M1539 293 30 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=136120 $D=0
M1540 294 30 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=140750 $D=0
M1541 295 30 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=145380 $D=0
M1542 163 31 296 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=136120 $D=0
M1543 167 31 297 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=140750 $D=0
M1544 168 31 298 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=145380 $D=0
M1545 299 32 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=136120 $D=0
M1546 300 32 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=140750 $D=0
M1547 301 32 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=145380 $D=0
M1548 302 296 227 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=136120 $D=0
M1549 303 297 228 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=140750 $D=0
M1550 304 298 229 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=145380 $D=0
M1551 163 302 957 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=136120 $D=0
M1552 167 303 958 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=140750 $D=0
M1553 168 304 959 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=145380 $D=0
M1554 305 957 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=136120 $D=0
M1555 306 958 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=140750 $D=0
M1556 307 959 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=145380 $D=0
M1557 302 31 305 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=136120 $D=0
M1558 303 31 306 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=140750 $D=0
M1559 304 31 307 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=145380 $D=0
M1560 305 299 242 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=136120 $D=0
M1561 306 300 243 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=140750 $D=0
M1562 307 301 244 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=145380 $D=0
M1563 248 308 305 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=136120 $D=0
M1564 249 309 306 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=140750 $D=0
M1565 250 310 307 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=145380 $D=0
M1566 308 33 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=136120 $D=0
M1567 309 33 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=140750 $D=0
M1568 310 33 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=145380 $D=0
M1569 163 34 311 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=136120 $D=0
M1570 167 34 312 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=140750 $D=0
M1571 168 34 313 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=145380 $D=0
M1572 314 35 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=136120 $D=0
M1573 315 35 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=140750 $D=0
M1574 316 35 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=145380 $D=0
M1575 317 311 227 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=136120 $D=0
M1576 318 312 228 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=140750 $D=0
M1577 319 313 229 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=145380 $D=0
M1578 163 317 960 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=136120 $D=0
M1579 167 318 961 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=140750 $D=0
M1580 168 319 962 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=145380 $D=0
M1581 320 960 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=136120 $D=0
M1582 321 961 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=140750 $D=0
M1583 322 962 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=145380 $D=0
M1584 317 34 320 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=136120 $D=0
M1585 318 34 321 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=140750 $D=0
M1586 319 34 322 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=145380 $D=0
M1587 320 314 242 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=136120 $D=0
M1588 321 315 243 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=140750 $D=0
M1589 322 316 244 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=145380 $D=0
M1590 248 323 320 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=136120 $D=0
M1591 249 324 321 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=140750 $D=0
M1592 250 325 322 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=145380 $D=0
M1593 323 36 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=136120 $D=0
M1594 324 36 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=140750 $D=0
M1595 325 36 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=145380 $D=0
M1596 163 37 326 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=136120 $D=0
M1597 167 37 327 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=140750 $D=0
M1598 168 37 328 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=145380 $D=0
M1599 329 38 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=136120 $D=0
M1600 330 38 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=140750 $D=0
M1601 331 38 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=145380 $D=0
M1602 332 326 227 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=136120 $D=0
M1603 333 327 228 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=140750 $D=0
M1604 334 328 229 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=145380 $D=0
M1605 163 332 963 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=136120 $D=0
M1606 167 333 964 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=140750 $D=0
M1607 168 334 965 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=145380 $D=0
M1608 335 963 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=136120 $D=0
M1609 336 964 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=140750 $D=0
M1610 337 965 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=145380 $D=0
M1611 332 37 335 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=136120 $D=0
M1612 333 37 336 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=140750 $D=0
M1613 334 37 337 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=145380 $D=0
M1614 335 329 242 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=136120 $D=0
M1615 336 330 243 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=140750 $D=0
M1616 337 331 244 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=145380 $D=0
M1617 248 338 335 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=136120 $D=0
M1618 249 339 336 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=140750 $D=0
M1619 250 340 337 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=145380 $D=0
M1620 338 39 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=136120 $D=0
M1621 339 39 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=140750 $D=0
M1622 340 39 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=145380 $D=0
M1623 163 40 341 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=136120 $D=0
M1624 167 40 342 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=140750 $D=0
M1625 168 40 343 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=145380 $D=0
M1626 344 41 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=136120 $D=0
M1627 345 41 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=140750 $D=0
M1628 346 41 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=145380 $D=0
M1629 347 341 227 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=136120 $D=0
M1630 348 342 228 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=140750 $D=0
M1631 349 343 229 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=145380 $D=0
M1632 163 347 966 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=136120 $D=0
M1633 167 348 967 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=140750 $D=0
M1634 168 349 968 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=145380 $D=0
M1635 350 966 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=136120 $D=0
M1636 351 967 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=140750 $D=0
M1637 352 968 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=145380 $D=0
M1638 347 40 350 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=136120 $D=0
M1639 348 40 351 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=140750 $D=0
M1640 349 40 352 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=145380 $D=0
M1641 350 344 242 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=136120 $D=0
M1642 351 345 243 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=140750 $D=0
M1643 352 346 244 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=145380 $D=0
M1644 248 353 350 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=136120 $D=0
M1645 249 354 351 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=140750 $D=0
M1646 250 355 352 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=145380 $D=0
M1647 353 42 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=136120 $D=0
M1648 354 42 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=140750 $D=0
M1649 355 42 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=145380 $D=0
M1650 163 43 356 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=136120 $D=0
M1651 167 43 357 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=140750 $D=0
M1652 168 43 358 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=145380 $D=0
M1653 359 44 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=136120 $D=0
M1654 360 44 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=140750 $D=0
M1655 361 44 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=145380 $D=0
M1656 362 356 227 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=136120 $D=0
M1657 363 357 228 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=140750 $D=0
M1658 364 358 229 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=145380 $D=0
M1659 163 362 969 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=136120 $D=0
M1660 167 363 970 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=140750 $D=0
M1661 168 364 971 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=145380 $D=0
M1662 365 969 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=136120 $D=0
M1663 366 970 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=140750 $D=0
M1664 367 971 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=145380 $D=0
M1665 362 43 365 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=136120 $D=0
M1666 363 43 366 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=140750 $D=0
M1667 364 43 367 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=145380 $D=0
M1668 365 359 242 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=136120 $D=0
M1669 366 360 243 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=140750 $D=0
M1670 367 361 244 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=145380 $D=0
M1671 248 368 365 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=136120 $D=0
M1672 249 369 366 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=140750 $D=0
M1673 250 370 367 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=145380 $D=0
M1674 368 45 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=136120 $D=0
M1675 369 45 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=140750 $D=0
M1676 370 45 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=145380 $D=0
M1677 163 46 371 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=136120 $D=0
M1678 167 46 372 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=140750 $D=0
M1679 168 46 373 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=145380 $D=0
M1680 374 47 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=136120 $D=0
M1681 375 47 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=140750 $D=0
M1682 376 47 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=145380 $D=0
M1683 377 371 227 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=136120 $D=0
M1684 378 372 228 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=140750 $D=0
M1685 379 373 229 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=145380 $D=0
M1686 163 377 972 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=136120 $D=0
M1687 167 378 973 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=140750 $D=0
M1688 168 379 974 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=145380 $D=0
M1689 380 972 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=136120 $D=0
M1690 381 973 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=140750 $D=0
M1691 382 974 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=145380 $D=0
M1692 377 46 380 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=136120 $D=0
M1693 378 46 381 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=140750 $D=0
M1694 379 46 382 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=145380 $D=0
M1695 380 374 242 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=136120 $D=0
M1696 381 375 243 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=140750 $D=0
M1697 382 376 244 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=145380 $D=0
M1698 248 383 380 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=136120 $D=0
M1699 249 384 381 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=140750 $D=0
M1700 250 385 382 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=145380 $D=0
M1701 383 48 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=136120 $D=0
M1702 384 48 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=140750 $D=0
M1703 385 48 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=145380 $D=0
M1704 163 49 386 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=136120 $D=0
M1705 167 49 387 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=140750 $D=0
M1706 168 49 388 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=145380 $D=0
M1707 389 50 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=136120 $D=0
M1708 390 50 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=140750 $D=0
M1709 391 50 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=145380 $D=0
M1710 392 386 227 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=136120 $D=0
M1711 393 387 228 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=140750 $D=0
M1712 394 388 229 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=145380 $D=0
M1713 163 392 975 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=136120 $D=0
M1714 167 393 976 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=140750 $D=0
M1715 168 394 977 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=145380 $D=0
M1716 395 975 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=136120 $D=0
M1717 396 976 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=140750 $D=0
M1718 397 977 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=145380 $D=0
M1719 392 49 395 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=136120 $D=0
M1720 393 49 396 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=140750 $D=0
M1721 394 49 397 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=145380 $D=0
M1722 395 389 242 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=136120 $D=0
M1723 396 390 243 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=140750 $D=0
M1724 397 391 244 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=145380 $D=0
M1725 248 398 395 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=136120 $D=0
M1726 249 399 396 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=140750 $D=0
M1727 250 400 397 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=145380 $D=0
M1728 398 51 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=136120 $D=0
M1729 399 51 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=140750 $D=0
M1730 400 51 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=145380 $D=0
M1731 163 52 401 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=136120 $D=0
M1732 167 52 402 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=140750 $D=0
M1733 168 52 403 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=145380 $D=0
M1734 404 53 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=136120 $D=0
M1735 405 53 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=140750 $D=0
M1736 406 53 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=145380 $D=0
M1737 407 401 227 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=136120 $D=0
M1738 408 402 228 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=140750 $D=0
M1739 409 403 229 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=145380 $D=0
M1740 163 407 978 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=136120 $D=0
M1741 167 408 979 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=140750 $D=0
M1742 168 409 980 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=145380 $D=0
M1743 410 978 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=136120 $D=0
M1744 411 979 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=140750 $D=0
M1745 412 980 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=145380 $D=0
M1746 407 52 410 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=136120 $D=0
M1747 408 52 411 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=140750 $D=0
M1748 409 52 412 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=145380 $D=0
M1749 410 404 242 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=136120 $D=0
M1750 411 405 243 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=140750 $D=0
M1751 412 406 244 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=145380 $D=0
M1752 248 413 410 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=136120 $D=0
M1753 249 414 411 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=140750 $D=0
M1754 250 415 412 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=145380 $D=0
M1755 413 54 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=136120 $D=0
M1756 414 54 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=140750 $D=0
M1757 415 54 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=145380 $D=0
M1758 163 55 416 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=136120 $D=0
M1759 167 55 417 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=140750 $D=0
M1760 168 55 418 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=145380 $D=0
M1761 419 56 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=136120 $D=0
M1762 420 56 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=140750 $D=0
M1763 421 56 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=145380 $D=0
M1764 422 416 227 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=136120 $D=0
M1765 423 417 228 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=140750 $D=0
M1766 424 418 229 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=145380 $D=0
M1767 163 422 981 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=136120 $D=0
M1768 167 423 982 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=140750 $D=0
M1769 168 424 983 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=145380 $D=0
M1770 425 981 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=136120 $D=0
M1771 426 982 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=140750 $D=0
M1772 427 983 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=145380 $D=0
M1773 422 55 425 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=136120 $D=0
M1774 423 55 426 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=140750 $D=0
M1775 424 55 427 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=145380 $D=0
M1776 425 419 242 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=136120 $D=0
M1777 426 420 243 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=140750 $D=0
M1778 427 421 244 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=145380 $D=0
M1779 248 428 425 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=136120 $D=0
M1780 249 429 426 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=140750 $D=0
M1781 250 430 427 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=145380 $D=0
M1782 428 57 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=136120 $D=0
M1783 429 57 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=140750 $D=0
M1784 430 57 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=145380 $D=0
M1785 163 58 431 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=136120 $D=0
M1786 167 58 432 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=140750 $D=0
M1787 168 58 433 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=145380 $D=0
M1788 434 59 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=136120 $D=0
M1789 435 59 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=140750 $D=0
M1790 436 59 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=145380 $D=0
M1791 437 431 227 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=136120 $D=0
M1792 438 432 228 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=140750 $D=0
M1793 439 433 229 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=145380 $D=0
M1794 163 437 984 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=136120 $D=0
M1795 167 438 985 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=140750 $D=0
M1796 168 439 986 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=145380 $D=0
M1797 440 984 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=136120 $D=0
M1798 441 985 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=140750 $D=0
M1799 442 986 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=145380 $D=0
M1800 437 58 440 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=136120 $D=0
M1801 438 58 441 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=140750 $D=0
M1802 439 58 442 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=145380 $D=0
M1803 440 434 242 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=136120 $D=0
M1804 441 435 243 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=140750 $D=0
M1805 442 436 244 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=145380 $D=0
M1806 248 443 440 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=136120 $D=0
M1807 249 444 441 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=140750 $D=0
M1808 250 445 442 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=145380 $D=0
M1809 443 60 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=136120 $D=0
M1810 444 60 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=140750 $D=0
M1811 445 60 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=145380 $D=0
M1812 163 61 446 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=136120 $D=0
M1813 167 61 447 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=140750 $D=0
M1814 168 61 448 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=145380 $D=0
M1815 449 62 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=136120 $D=0
M1816 450 62 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=140750 $D=0
M1817 451 62 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=145380 $D=0
M1818 452 446 227 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=136120 $D=0
M1819 453 447 228 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=140750 $D=0
M1820 454 448 229 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=145380 $D=0
M1821 163 452 987 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=136120 $D=0
M1822 167 453 988 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=140750 $D=0
M1823 168 454 989 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=145380 $D=0
M1824 455 987 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=136120 $D=0
M1825 456 988 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=140750 $D=0
M1826 457 989 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=145380 $D=0
M1827 452 61 455 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=136120 $D=0
M1828 453 61 456 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=140750 $D=0
M1829 454 61 457 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=145380 $D=0
M1830 455 449 242 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=136120 $D=0
M1831 456 450 243 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=140750 $D=0
M1832 457 451 244 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=145380 $D=0
M1833 248 458 455 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=136120 $D=0
M1834 249 459 456 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=140750 $D=0
M1835 250 460 457 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=145380 $D=0
M1836 458 63 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=136120 $D=0
M1837 459 63 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=140750 $D=0
M1838 460 63 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=145380 $D=0
M1839 163 64 461 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=136120 $D=0
M1840 167 64 462 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=140750 $D=0
M1841 168 64 463 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=145380 $D=0
M1842 464 65 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=136120 $D=0
M1843 465 65 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=140750 $D=0
M1844 466 65 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=145380 $D=0
M1845 467 461 227 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=136120 $D=0
M1846 468 462 228 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=140750 $D=0
M1847 469 463 229 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=145380 $D=0
M1848 163 467 990 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=136120 $D=0
M1849 167 468 991 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=140750 $D=0
M1850 168 469 992 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=145380 $D=0
M1851 470 990 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=136120 $D=0
M1852 471 991 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=140750 $D=0
M1853 472 992 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=145380 $D=0
M1854 467 64 470 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=136120 $D=0
M1855 468 64 471 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=140750 $D=0
M1856 469 64 472 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=145380 $D=0
M1857 470 464 242 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=136120 $D=0
M1858 471 465 243 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=140750 $D=0
M1859 472 466 244 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=145380 $D=0
M1860 248 473 470 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=136120 $D=0
M1861 249 474 471 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=140750 $D=0
M1862 250 475 472 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=145380 $D=0
M1863 473 66 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=136120 $D=0
M1864 474 66 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=140750 $D=0
M1865 475 66 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=145380 $D=0
M1866 163 67 476 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=136120 $D=0
M1867 167 67 477 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=140750 $D=0
M1868 168 67 478 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=145380 $D=0
M1869 479 68 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=136120 $D=0
M1870 480 68 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=140750 $D=0
M1871 481 68 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=145380 $D=0
M1872 482 476 227 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=136120 $D=0
M1873 483 477 228 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=140750 $D=0
M1874 484 478 229 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=145380 $D=0
M1875 163 482 993 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=136120 $D=0
M1876 167 483 994 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=140750 $D=0
M1877 168 484 995 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=145380 $D=0
M1878 485 993 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=136120 $D=0
M1879 486 994 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=140750 $D=0
M1880 487 995 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=145380 $D=0
M1881 482 67 485 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=136120 $D=0
M1882 483 67 486 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=140750 $D=0
M1883 484 67 487 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=145380 $D=0
M1884 485 479 242 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=136120 $D=0
M1885 486 480 243 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=140750 $D=0
M1886 487 481 244 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=145380 $D=0
M1887 248 488 485 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=136120 $D=0
M1888 249 489 486 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=140750 $D=0
M1889 250 490 487 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=145380 $D=0
M1890 488 69 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=136120 $D=0
M1891 489 69 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=140750 $D=0
M1892 490 69 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=145380 $D=0
M1893 163 70 491 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=136120 $D=0
M1894 167 70 492 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=140750 $D=0
M1895 168 70 493 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=145380 $D=0
M1896 494 71 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=136120 $D=0
M1897 495 71 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=140750 $D=0
M1898 496 71 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=145380 $D=0
M1899 497 491 227 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=136120 $D=0
M1900 498 492 228 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=140750 $D=0
M1901 499 493 229 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=145380 $D=0
M1902 163 497 996 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=136120 $D=0
M1903 167 498 997 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=140750 $D=0
M1904 168 499 998 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=145380 $D=0
M1905 500 996 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=136120 $D=0
M1906 501 997 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=140750 $D=0
M1907 502 998 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=145380 $D=0
M1908 497 70 500 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=136120 $D=0
M1909 498 70 501 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=140750 $D=0
M1910 499 70 502 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=145380 $D=0
M1911 500 494 242 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=136120 $D=0
M1912 501 495 243 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=140750 $D=0
M1913 502 496 244 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=145380 $D=0
M1914 248 503 500 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=136120 $D=0
M1915 249 504 501 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=140750 $D=0
M1916 250 505 502 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=145380 $D=0
M1917 503 72 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=136120 $D=0
M1918 504 72 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=140750 $D=0
M1919 505 72 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=145380 $D=0
M1920 163 73 506 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=136120 $D=0
M1921 167 73 507 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=140750 $D=0
M1922 168 73 508 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=145380 $D=0
M1923 509 74 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=136120 $D=0
M1924 510 74 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=140750 $D=0
M1925 511 74 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=145380 $D=0
M1926 512 506 227 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=136120 $D=0
M1927 513 507 228 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=140750 $D=0
M1928 514 508 229 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=145380 $D=0
M1929 163 512 999 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=136120 $D=0
M1930 167 513 1000 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=140750 $D=0
M1931 168 514 1001 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=145380 $D=0
M1932 515 999 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=136120 $D=0
M1933 516 1000 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=140750 $D=0
M1934 517 1001 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=145380 $D=0
M1935 512 73 515 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=136120 $D=0
M1936 513 73 516 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=140750 $D=0
M1937 514 73 517 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=145380 $D=0
M1938 515 509 242 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=136120 $D=0
M1939 516 510 243 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=140750 $D=0
M1940 517 511 244 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=145380 $D=0
M1941 248 518 515 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=136120 $D=0
M1942 249 519 516 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=140750 $D=0
M1943 250 520 517 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=145380 $D=0
M1944 518 75 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=136120 $D=0
M1945 519 75 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=140750 $D=0
M1946 520 75 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=145380 $D=0
M1947 163 76 521 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=136120 $D=0
M1948 167 76 522 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=140750 $D=0
M1949 168 76 523 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=145380 $D=0
M1950 524 77 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=136120 $D=0
M1951 525 77 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=140750 $D=0
M1952 526 77 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=145380 $D=0
M1953 527 521 227 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=136120 $D=0
M1954 528 522 228 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=140750 $D=0
M1955 529 523 229 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=145380 $D=0
M1956 163 527 1002 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=136120 $D=0
M1957 167 528 1003 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=140750 $D=0
M1958 168 529 1004 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=145380 $D=0
M1959 530 1002 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=136120 $D=0
M1960 531 1003 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=140750 $D=0
M1961 532 1004 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=145380 $D=0
M1962 527 76 530 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=136120 $D=0
M1963 528 76 531 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=140750 $D=0
M1964 529 76 532 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=145380 $D=0
M1965 530 524 242 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=136120 $D=0
M1966 531 525 243 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=140750 $D=0
M1967 532 526 244 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=145380 $D=0
M1968 248 533 530 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=136120 $D=0
M1969 249 534 531 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=140750 $D=0
M1970 250 535 532 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=145380 $D=0
M1971 533 78 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=136120 $D=0
M1972 534 78 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=140750 $D=0
M1973 535 78 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=145380 $D=0
M1974 163 79 536 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=136120 $D=0
M1975 167 79 537 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=140750 $D=0
M1976 168 79 538 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=145380 $D=0
M1977 539 80 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=136120 $D=0
M1978 540 80 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=140750 $D=0
M1979 541 80 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=145380 $D=0
M1980 542 536 227 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=136120 $D=0
M1981 543 537 228 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=140750 $D=0
M1982 544 538 229 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=145380 $D=0
M1983 163 542 1005 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=136120 $D=0
M1984 167 543 1006 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=140750 $D=0
M1985 168 544 1007 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=145380 $D=0
M1986 545 1005 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=136120 $D=0
M1987 546 1006 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=140750 $D=0
M1988 547 1007 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=145380 $D=0
M1989 542 79 545 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=136120 $D=0
M1990 543 79 546 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=140750 $D=0
M1991 544 79 547 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=145380 $D=0
M1992 545 539 242 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=136120 $D=0
M1993 546 540 243 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=140750 $D=0
M1994 547 541 244 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=145380 $D=0
M1995 248 548 545 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=136120 $D=0
M1996 249 549 546 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=140750 $D=0
M1997 250 550 547 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=145380 $D=0
M1998 548 81 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=136120 $D=0
M1999 549 81 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=140750 $D=0
M2000 550 81 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=145380 $D=0
M2001 163 82 551 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=136120 $D=0
M2002 167 82 552 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=140750 $D=0
M2003 168 82 553 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=145380 $D=0
M2004 554 83 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=136120 $D=0
M2005 555 83 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=140750 $D=0
M2006 556 83 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=145380 $D=0
M2007 557 551 227 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=136120 $D=0
M2008 558 552 228 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=140750 $D=0
M2009 559 553 229 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=145380 $D=0
M2010 163 557 1008 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=136120 $D=0
M2011 167 558 1009 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=140750 $D=0
M2012 168 559 1010 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=145380 $D=0
M2013 560 1008 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=136120 $D=0
M2014 561 1009 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=140750 $D=0
M2015 562 1010 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=145380 $D=0
M2016 557 82 560 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=136120 $D=0
M2017 558 82 561 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=140750 $D=0
M2018 559 82 562 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=145380 $D=0
M2019 560 554 242 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=136120 $D=0
M2020 561 555 243 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=140750 $D=0
M2021 562 556 244 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=145380 $D=0
M2022 248 563 560 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=136120 $D=0
M2023 249 564 561 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=140750 $D=0
M2024 250 565 562 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=145380 $D=0
M2025 563 84 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=136120 $D=0
M2026 564 84 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=140750 $D=0
M2027 565 84 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=145380 $D=0
M2028 163 85 566 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=136120 $D=0
M2029 167 85 567 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=140750 $D=0
M2030 168 85 568 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=145380 $D=0
M2031 569 86 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=136120 $D=0
M2032 570 86 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=140750 $D=0
M2033 571 86 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=145380 $D=0
M2034 572 566 227 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=136120 $D=0
M2035 573 567 228 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=140750 $D=0
M2036 574 568 229 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=145380 $D=0
M2037 163 572 1011 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=136120 $D=0
M2038 167 573 1012 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=140750 $D=0
M2039 168 574 1013 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=145380 $D=0
M2040 575 1011 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=136120 $D=0
M2041 576 1012 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=140750 $D=0
M2042 577 1013 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=145380 $D=0
M2043 572 85 575 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=136120 $D=0
M2044 573 85 576 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=140750 $D=0
M2045 574 85 577 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=145380 $D=0
M2046 575 569 242 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=136120 $D=0
M2047 576 570 243 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=140750 $D=0
M2048 577 571 244 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=145380 $D=0
M2049 248 578 575 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=136120 $D=0
M2050 249 579 576 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=140750 $D=0
M2051 250 580 577 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=145380 $D=0
M2052 578 87 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=136120 $D=0
M2053 579 87 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=140750 $D=0
M2054 580 87 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=145380 $D=0
M2055 163 88 581 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=136120 $D=0
M2056 167 88 582 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=140750 $D=0
M2057 168 88 583 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=145380 $D=0
M2058 584 89 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=136120 $D=0
M2059 585 89 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=140750 $D=0
M2060 586 89 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=145380 $D=0
M2061 587 581 227 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=136120 $D=0
M2062 588 582 228 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=140750 $D=0
M2063 589 583 229 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=145380 $D=0
M2064 163 587 1014 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=136120 $D=0
M2065 167 588 1015 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=140750 $D=0
M2066 168 589 1016 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=145380 $D=0
M2067 590 1014 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=136120 $D=0
M2068 591 1015 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=140750 $D=0
M2069 592 1016 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=145380 $D=0
M2070 587 88 590 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=136120 $D=0
M2071 588 88 591 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=140750 $D=0
M2072 589 88 592 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=145380 $D=0
M2073 590 584 242 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=136120 $D=0
M2074 591 585 243 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=140750 $D=0
M2075 592 586 244 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=145380 $D=0
M2076 248 593 590 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=136120 $D=0
M2077 249 594 591 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=140750 $D=0
M2078 250 595 592 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=145380 $D=0
M2079 593 90 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=136120 $D=0
M2080 594 90 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=140750 $D=0
M2081 595 90 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=145380 $D=0
M2082 163 91 596 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=136120 $D=0
M2083 167 91 597 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=140750 $D=0
M2084 168 91 598 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=145380 $D=0
M2085 599 92 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=136120 $D=0
M2086 600 92 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=140750 $D=0
M2087 601 92 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=145380 $D=0
M2088 602 596 227 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=136120 $D=0
M2089 603 597 228 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=140750 $D=0
M2090 604 598 229 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=145380 $D=0
M2091 163 602 1017 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=136120 $D=0
M2092 167 603 1018 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=140750 $D=0
M2093 168 604 1019 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=145380 $D=0
M2094 605 1017 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=136120 $D=0
M2095 606 1018 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=140750 $D=0
M2096 607 1019 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=145380 $D=0
M2097 602 91 605 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=136120 $D=0
M2098 603 91 606 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=140750 $D=0
M2099 604 91 607 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=145380 $D=0
M2100 605 599 242 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=136120 $D=0
M2101 606 600 243 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=140750 $D=0
M2102 607 601 244 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=145380 $D=0
M2103 248 608 605 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=136120 $D=0
M2104 249 609 606 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=140750 $D=0
M2105 250 610 607 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=145380 $D=0
M2106 608 93 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=136120 $D=0
M2107 609 93 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=140750 $D=0
M2108 610 93 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=145380 $D=0
M2109 163 94 611 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=136120 $D=0
M2110 167 94 612 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=140750 $D=0
M2111 168 94 613 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=145380 $D=0
M2112 614 95 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=136120 $D=0
M2113 615 95 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=140750 $D=0
M2114 616 95 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=145380 $D=0
M2115 617 611 227 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=136120 $D=0
M2116 618 612 228 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=140750 $D=0
M2117 619 613 229 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=145380 $D=0
M2118 163 617 1020 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=136120 $D=0
M2119 167 618 1021 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=140750 $D=0
M2120 168 619 1022 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=145380 $D=0
M2121 620 1020 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=136120 $D=0
M2122 621 1021 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=140750 $D=0
M2123 622 1022 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=145380 $D=0
M2124 617 94 620 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=136120 $D=0
M2125 618 94 621 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=140750 $D=0
M2126 619 94 622 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=145380 $D=0
M2127 620 614 242 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=136120 $D=0
M2128 621 615 243 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=140750 $D=0
M2129 622 616 244 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=145380 $D=0
M2130 248 623 620 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=136120 $D=0
M2131 249 624 621 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=140750 $D=0
M2132 250 625 622 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=145380 $D=0
M2133 623 96 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=136120 $D=0
M2134 624 96 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=140750 $D=0
M2135 625 96 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=145380 $D=0
M2136 163 97 626 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=136120 $D=0
M2137 167 97 627 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=140750 $D=0
M2138 168 97 628 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=145380 $D=0
M2139 629 98 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=136120 $D=0
M2140 630 98 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=140750 $D=0
M2141 631 98 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=145380 $D=0
M2142 632 626 227 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=136120 $D=0
M2143 633 627 228 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=140750 $D=0
M2144 634 628 229 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=145380 $D=0
M2145 163 632 1023 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=136120 $D=0
M2146 167 633 1024 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=140750 $D=0
M2147 168 634 1025 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=145380 $D=0
M2148 635 1023 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=136120 $D=0
M2149 636 1024 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=140750 $D=0
M2150 637 1025 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=145380 $D=0
M2151 632 97 635 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=136120 $D=0
M2152 633 97 636 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=140750 $D=0
M2153 634 97 637 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=145380 $D=0
M2154 635 629 242 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=136120 $D=0
M2155 636 630 243 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=140750 $D=0
M2156 637 631 244 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=145380 $D=0
M2157 248 638 635 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=136120 $D=0
M2158 249 639 636 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=140750 $D=0
M2159 250 640 637 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=145380 $D=0
M2160 638 99 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=136120 $D=0
M2161 639 99 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=140750 $D=0
M2162 640 99 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=145380 $D=0
M2163 163 100 641 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=136120 $D=0
M2164 167 100 642 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=140750 $D=0
M2165 168 100 643 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=145380 $D=0
M2166 644 101 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=136120 $D=0
M2167 645 101 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=140750 $D=0
M2168 646 101 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=145380 $D=0
M2169 647 641 227 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=136120 $D=0
M2170 648 642 228 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=140750 $D=0
M2171 649 643 229 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=145380 $D=0
M2172 163 647 1026 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=136120 $D=0
M2173 167 648 1027 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=140750 $D=0
M2174 168 649 1028 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=145380 $D=0
M2175 650 1026 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=136120 $D=0
M2176 651 1027 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=140750 $D=0
M2177 652 1028 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=145380 $D=0
M2178 647 100 650 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=136120 $D=0
M2179 648 100 651 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=140750 $D=0
M2180 649 100 652 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=145380 $D=0
M2181 650 644 242 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=136120 $D=0
M2182 651 645 243 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=140750 $D=0
M2183 652 646 244 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=145380 $D=0
M2184 248 653 650 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=136120 $D=0
M2185 249 654 651 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=140750 $D=0
M2186 250 655 652 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=145380 $D=0
M2187 653 102 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=136120 $D=0
M2188 654 102 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=140750 $D=0
M2189 655 102 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=145380 $D=0
M2190 163 103 656 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=136120 $D=0
M2191 167 103 657 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=140750 $D=0
M2192 168 103 658 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=145380 $D=0
M2193 659 104 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=136120 $D=0
M2194 660 104 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=140750 $D=0
M2195 661 104 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=145380 $D=0
M2196 662 656 227 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=136120 $D=0
M2197 663 657 228 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=140750 $D=0
M2198 664 658 229 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=145380 $D=0
M2199 163 662 1029 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=136120 $D=0
M2200 167 663 1030 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=140750 $D=0
M2201 168 664 1031 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=145380 $D=0
M2202 665 1029 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=136120 $D=0
M2203 666 1030 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=140750 $D=0
M2204 667 1031 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=145380 $D=0
M2205 662 103 665 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=136120 $D=0
M2206 663 103 666 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=140750 $D=0
M2207 664 103 667 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=145380 $D=0
M2208 665 659 242 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=136120 $D=0
M2209 666 660 243 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=140750 $D=0
M2210 667 661 244 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=145380 $D=0
M2211 248 668 665 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=136120 $D=0
M2212 249 669 666 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=140750 $D=0
M2213 250 670 667 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=145380 $D=0
M2214 668 105 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=136120 $D=0
M2215 669 105 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=140750 $D=0
M2216 670 105 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=145380 $D=0
M2217 163 106 671 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=136120 $D=0
M2218 167 106 672 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=140750 $D=0
M2219 168 106 673 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=145380 $D=0
M2220 674 107 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=136120 $D=0
M2221 675 107 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=140750 $D=0
M2222 676 107 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=145380 $D=0
M2223 677 671 227 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=136120 $D=0
M2224 678 672 228 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=140750 $D=0
M2225 679 673 229 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=145380 $D=0
M2226 163 677 1032 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=136120 $D=0
M2227 167 678 1033 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=140750 $D=0
M2228 168 679 1034 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=145380 $D=0
M2229 680 1032 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=136120 $D=0
M2230 681 1033 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=140750 $D=0
M2231 682 1034 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=145380 $D=0
M2232 677 106 680 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=136120 $D=0
M2233 678 106 681 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=140750 $D=0
M2234 679 106 682 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=145380 $D=0
M2235 680 674 242 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=136120 $D=0
M2236 681 675 243 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=140750 $D=0
M2237 682 676 244 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=145380 $D=0
M2238 248 683 680 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=136120 $D=0
M2239 249 684 681 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=140750 $D=0
M2240 250 685 682 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=145380 $D=0
M2241 683 108 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=136120 $D=0
M2242 684 108 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=140750 $D=0
M2243 685 108 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=145380 $D=0
M2244 163 109 686 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=136120 $D=0
M2245 167 109 687 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=140750 $D=0
M2246 168 109 688 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=145380 $D=0
M2247 689 110 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=136120 $D=0
M2248 690 110 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=140750 $D=0
M2249 691 110 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=145380 $D=0
M2250 692 686 227 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=136120 $D=0
M2251 693 687 228 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=140750 $D=0
M2252 694 688 229 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=145380 $D=0
M2253 163 692 1035 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=136120 $D=0
M2254 167 693 1036 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=140750 $D=0
M2255 168 694 1037 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=145380 $D=0
M2256 695 1035 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=136120 $D=0
M2257 696 1036 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=140750 $D=0
M2258 697 1037 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=145380 $D=0
M2259 692 109 695 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=136120 $D=0
M2260 693 109 696 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=140750 $D=0
M2261 694 109 697 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=145380 $D=0
M2262 695 689 242 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=136120 $D=0
M2263 696 690 243 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=140750 $D=0
M2264 697 691 244 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=145380 $D=0
M2265 248 698 695 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=136120 $D=0
M2266 249 699 696 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=140750 $D=0
M2267 250 700 697 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=145380 $D=0
M2268 698 111 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=136120 $D=0
M2269 699 111 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=140750 $D=0
M2270 700 111 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=145380 $D=0
M2271 163 112 701 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=136120 $D=0
M2272 167 112 702 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=140750 $D=0
M2273 168 112 703 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=145380 $D=0
M2274 704 113 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=136120 $D=0
M2275 705 113 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=140750 $D=0
M2276 706 113 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=145380 $D=0
M2277 8 704 242 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=136120 $D=0
M2278 9 705 243 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=140750 $D=0
M2279 136 706 244 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=145380 $D=0
M2280 248 701 8 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=136120 $D=0
M2281 249 702 9 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=140750 $D=0
M2282 250 703 136 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=145380 $D=0
M2283 163 710 707 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=136120 $D=0
M2284 167 711 708 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=140750 $D=0
M2285 168 712 709 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=145380 $D=0
M2286 710 114 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=136120 $D=0
M2287 711 114 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=140750 $D=0
M2288 712 114 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=145380 $D=0
M2289 1038 242 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=136120 $D=0
M2290 1039 243 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=140750 $D=0
M2291 1040 244 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=145380 $D=0
M2292 713 710 1038 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=136120 $D=0
M2293 714 711 1039 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=140750 $D=0
M2294 715 712 1040 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=145380 $D=0
M2295 163 713 716 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=136120 $D=0
M2296 167 714 717 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=140750 $D=0
M2297 168 715 718 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=145380 $D=0
M2298 1041 716 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=136120 $D=0
M2299 1042 717 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=140750 $D=0
M2300 1043 718 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=145380 $D=0
M2301 713 707 1041 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=136120 $D=0
M2302 714 708 1042 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=140750 $D=0
M2303 715 709 1043 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=145380 $D=0
M2304 163 722 719 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=136120 $D=0
M2305 167 723 720 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=140750 $D=0
M2306 168 724 721 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=145380 $D=0
M2307 722 114 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=136120 $D=0
M2308 723 114 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=140750 $D=0
M2309 724 114 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=145380 $D=0
M2310 1044 248 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=136120 $D=0
M2311 1045 249 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=140750 $D=0
M2312 1046 250 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=145380 $D=0
M2313 725 722 1044 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=136120 $D=0
M2314 726 723 1045 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=140750 $D=0
M2315 727 724 1046 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=145380 $D=0
M2316 163 725 115 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=136120 $D=0
M2317 167 726 116 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=140750 $D=0
M2318 168 727 117 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=145380 $D=0
M2319 1047 115 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=136120 $D=0
M2320 1048 116 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=140750 $D=0
M2321 1049 117 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=145380 $D=0
M2322 725 719 1047 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=136120 $D=0
M2323 726 720 1048 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=140750 $D=0
M2324 727 721 1049 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=145380 $D=0
M2325 728 118 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=136120 $D=0
M2326 729 118 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=140750 $D=0
M2327 730 118 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=145380 $D=0
M2328 731 118 716 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=136120 $D=0
M2329 732 118 717 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=140750 $D=0
M2330 733 118 718 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=145380 $D=0
M2331 119 728 731 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=136120 $D=0
M2332 120 729 732 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=140750 $D=0
M2333 121 730 733 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=145380 $D=0
M2334 734 122 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=136120 $D=0
M2335 735 122 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=140750 $D=0
M2336 736 122 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=145380 $D=0
M2337 737 122 115 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=136120 $D=0
M2338 738 122 116 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=140750 $D=0
M2339 739 122 117 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=145380 $D=0
M2340 1050 734 737 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=136120 $D=0
M2341 1051 735 738 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=140750 $D=0
M2342 1052 736 739 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=145380 $D=0
M2343 163 115 1050 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=136120 $D=0
M2344 167 116 1051 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=140750 $D=0
M2345 168 117 1052 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=145380 $D=0
M2346 740 123 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=136120 $D=0
M2347 741 123 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=140750 $D=0
M2348 742 123 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=145380 $D=0
M2349 124 123 737 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=136120 $D=0
M2350 125 123 738 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=140750 $D=0
M2351 126 123 739 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=145380 $D=0
M2352 11 740 124 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=136120 $D=0
M2353 12 741 125 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=140750 $D=0
M2354 13 742 126 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=145380 $D=0
M2355 745 743 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=136120 $D=0
M2356 746 744 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=140750 $D=0
M2357 747 127 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=145380 $D=0
M2358 163 751 748 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=136120 $D=0
M2359 167 752 749 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=140750 $D=0
M2360 168 753 750 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=145380 $D=0
M2361 754 731 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=136120 $D=0
M2362 755 732 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=140750 $D=0
M2363 756 733 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=145380 $D=0
M2364 751 731 743 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=136120 $D=0
M2365 752 732 744 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=140750 $D=0
M2366 753 733 127 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=145380 $D=0
M2367 745 754 751 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=136120 $D=0
M2368 746 755 752 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=140750 $D=0
M2369 747 756 753 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=145380 $D=0
M2370 757 748 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=136120 $D=0
M2371 758 749 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=140750 $D=0
M2372 759 750 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=145380 $D=0
M2373 128 748 124 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=136120 $D=0
M2374 743 749 125 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=140750 $D=0
M2375 744 750 126 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=145380 $D=0
M2376 731 757 128 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=136120 $D=0
M2377 732 758 743 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=140750 $D=0
M2378 733 759 744 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=145380 $D=0
M2379 760 128 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=136120 $D=0
M2380 761 743 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=140750 $D=0
M2381 762 744 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=145380 $D=0
M2382 763 748 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=136120 $D=0
M2383 764 749 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=140750 $D=0
M2384 765 750 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=145380 $D=0
M2385 766 748 760 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=136120 $D=0
M2386 767 749 761 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=140750 $D=0
M2387 768 750 762 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=145380 $D=0
M2388 124 763 766 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=136120 $D=0
M2389 125 764 767 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=140750 $D=0
M2390 126 765 768 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=145380 $D=0
M2391 1080 731 163 163 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=135760 $D=0
M2392 1081 732 167 167 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=140390 $D=0
M2393 1082 733 168 168 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=145020 $D=0
M2394 769 124 1080 163 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=135760 $D=0
M2395 770 125 1081 167 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=140390 $D=0
M2396 771 126 1082 168 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=145020 $D=0
M2397 772 766 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=136120 $D=0
M2398 773 767 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=140750 $D=0
M2399 774 768 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=145380 $D=0
M2400 775 731 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=136120 $D=0
M2401 776 732 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=140750 $D=0
M2402 777 733 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=145380 $D=0
M2403 163 124 775 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=136120 $D=0
M2404 167 125 776 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=140750 $D=0
M2405 168 126 777 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=145380 $D=0
M2406 778 731 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=136120 $D=0
M2407 779 732 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=140750 $D=0
M2408 780 733 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=145380 $D=0
M2409 163 124 778 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=136120 $D=0
M2410 167 125 779 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=140750 $D=0
M2411 168 126 780 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=145380 $D=0
M2412 1083 731 163 163 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=135940 $D=0
M2413 1084 732 167 167 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=140570 $D=0
M2414 1085 733 168 168 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=145200 $D=0
M2415 784 124 1083 163 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=135940 $D=0
M2416 785 125 1084 167 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=140570 $D=0
M2417 786 126 1085 168 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=145200 $D=0
M2418 163 778 784 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=136120 $D=0
M2419 167 779 785 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=140750 $D=0
M2420 168 780 786 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=145380 $D=0
M2421 787 132 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=136120 $D=0
M2422 788 132 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=140750 $D=0
M2423 789 132 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=145380 $D=0
M2424 790 132 769 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=136120 $D=0
M2425 791 132 770 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=140750 $D=0
M2426 792 132 771 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=145380 $D=0
M2427 775 787 790 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=136120 $D=0
M2428 776 788 791 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=140750 $D=0
M2429 777 789 792 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=145380 $D=0
M2430 793 132 772 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=136120 $D=0
M2431 794 132 773 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=140750 $D=0
M2432 795 132 774 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=145380 $D=0
M2433 784 787 793 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=136120 $D=0
M2434 785 788 794 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=140750 $D=0
M2435 786 789 795 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=145380 $D=0
M2436 796 133 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=136120 $D=0
M2437 797 133 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=140750 $D=0
M2438 798 133 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=145380 $D=0
M2439 799 133 793 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=136120 $D=0
M2440 800 133 794 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=140750 $D=0
M2441 801 133 795 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=145380 $D=0
M2442 790 796 799 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=136120 $D=0
M2443 791 797 800 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=140750 $D=0
M2444 792 798 801 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=145380 $D=0
M2445 14 799 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=136120 $D=0
M2446 15 800 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=140750 $D=0
M2447 16 801 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=145380 $D=0
M2448 802 134 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=136120 $D=0
M2449 803 134 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=140750 $D=0
M2450 804 134 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=145380 $D=0
M2451 805 134 125 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=136120 $D=0
M2452 806 134 135 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=140750 $D=0
M2453 807 134 136 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=145380 $D=0
M2454 137 802 805 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=136120 $D=0
M2455 124 803 806 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=140750 $D=0
M2456 125 804 807 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=145380 $D=0
M2457 808 134 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=136120 $D=0
M2458 809 134 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=140750 $D=0
M2459 810 134 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=145380 $D=0
M2460 817 134 138 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=136120 $D=0
M2461 818 134 9 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=140750 $D=0
M2462 819 134 136 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=145380 $D=0
M2463 139 808 817 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=136120 $D=0
M2464 140 809 818 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=140750 $D=0
M2465 141 810 819 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=145380 $D=0
M2466 820 134 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=136120 $D=0
M2467 821 134 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=140750 $D=0
M2468 822 134 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=145380 $D=0
M2469 823 134 8 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=136120 $D=0
M2470 824 134 9 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=140750 $D=0
M2471 825 134 136 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=145380 $D=0
M2472 142 820 823 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=136120 $D=0
M2473 143 821 824 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=140750 $D=0
M2474 144 822 825 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=145380 $D=0
M2475 826 134 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=136120 $D=0
M2476 827 134 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=140750 $D=0
M2477 828 134 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=145380 $D=0
M2478 829 134 8 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=136120 $D=0
M2479 830 134 9 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=140750 $D=0
M2480 831 134 136 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=145380 $D=0
M2481 145 826 829 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=136120 $D=0
M2482 146 827 830 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=140750 $D=0
M2483 147 828 831 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=145380 $D=0
M2484 832 134 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=136120 $D=0
M2485 833 134 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=140750 $D=0
M2486 834 134 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=145380 $D=0
M2487 835 134 8 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=136120 $D=0
M2488 836 134 9 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=140750 $D=0
M2489 837 134 136 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=145380 $D=0
M2490 148 832 835 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=136120 $D=0
M2491 149 833 836 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=140750 $D=0
M2492 144 834 837 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=145380 $D=0
M2493 163 731 1065 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=136120 $D=0
M2494 167 732 1066 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=140750 $D=0
M2495 168 733 1067 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=145380 $D=0
M2496 124 1065 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=136120 $D=0
M2497 125 1066 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=140750 $D=0
M2498 135 1067 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=145380 $D=0
M2499 838 126 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=136120 $D=0
M2500 839 126 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=140750 $D=0
M2501 840 126 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=145380 $D=0
M2502 141 126 124 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=136120 $D=0
M2503 150 126 125 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=140750 $D=0
M2504 138 126 135 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=145380 $D=0
M2505 805 838 141 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=136120 $D=0
M2506 806 839 150 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=140750 $D=0
M2507 807 840 138 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=145380 $D=0
M2508 841 125 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=136120 $D=0
M2509 842 125 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=140750 $D=0
M2510 843 125 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=145380 $D=0
M2511 131 125 141 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=136120 $D=0
M2512 130 125 150 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=140750 $D=0
M2513 129 125 138 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=145380 $D=0
M2514 817 841 131 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=136120 $D=0
M2515 818 842 130 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=140750 $D=0
M2516 819 843 129 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=145380 $D=0
M2517 844 124 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=136120 $D=0
M2518 845 124 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=140750 $D=0
M2519 846 124 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=145380 $D=0
M2520 151 124 131 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=136120 $D=0
M2521 152 124 130 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=140750 $D=0
M2522 153 124 129 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=145380 $D=0
M2523 823 844 151 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=136120 $D=0
M2524 824 845 152 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=140750 $D=0
M2525 825 846 153 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=145380 $D=0
M2526 847 154 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=136120 $D=0
M2527 848 154 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=140750 $D=0
M2528 849 154 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=145380 $D=0
M2529 155 154 151 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=136120 $D=0
M2530 156 154 152 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=140750 $D=0
M2531 157 154 153 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=145380 $D=0
M2532 829 847 155 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=136120 $D=0
M2533 830 848 156 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=140750 $D=0
M2534 831 849 157 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=145380 $D=0
M2535 850 158 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=136120 $D=0
M2536 851 158 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=140750 $D=0
M2537 852 158 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=145380 $D=0
M2538 206 158 155 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=136120 $D=0
M2539 207 158 156 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=140750 $D=0
M2540 208 158 157 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=145380 $D=0
M2541 835 850 206 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=136120 $D=0
M2542 836 851 207 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=140750 $D=0
M2543 837 852 208 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=145380 $D=0
M2544 853 159 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=136120 $D=0
M2545 854 159 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=140750 $D=0
M2546 855 159 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=145380 $D=0
M2547 856 159 115 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=136120 $D=0
M2548 857 159 116 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=140750 $D=0
M2549 858 159 117 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=145380 $D=0
M2550 11 853 856 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=136120 $D=0
M2551 12 854 857 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=140750 $D=0
M2552 13 855 858 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=145380 $D=0
M2553 859 716 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=136120 $D=0
M2554 860 717 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=140750 $D=0
M2555 861 718 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=145380 $D=0
M2556 163 856 859 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=136120 $D=0
M2557 167 857 860 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=140750 $D=0
M2558 168 858 861 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=145380 $D=0
M2559 1086 716 163 163 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=135940 $D=0
M2560 1087 717 167 167 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=140570 $D=0
M2561 1088 718 168 168 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=145200 $D=0
M2562 865 856 1086 163 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=135940 $D=0
M2563 866 857 1087 167 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=140570 $D=0
M2564 867 858 1088 168 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=145200 $D=0
M2565 163 859 865 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=136120 $D=0
M2566 167 860 866 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=140750 $D=0
M2567 168 861 867 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=145380 $D=0
M2568 1068 868 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=136120 $D=0
M2569 1069 869 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=140750 $D=0
M2570 1070 870 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=145380 $D=0
M2571 163 865 1068 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=136120 $D=0
M2572 167 866 1069 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=140750 $D=0
M2573 168 867 1070 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=145380 $D=0
M2574 869 1068 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=136120 $D=0
M2575 871 1069 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=140750 $D=0
M2576 160 1070 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=145380 $D=0
M2577 1089 716 163 163 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=135760 $D=0
M2578 1090 717 167 167 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=140390 $D=0
M2579 1091 718 168 168 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=145020 $D=0
M2580 872 875 1089 163 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=135760 $D=0
M2581 873 876 1090 167 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=140390 $D=0
M2582 874 877 1091 168 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=145020 $D=0
M2583 875 856 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=136120 $D=0
M2584 876 857 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=140750 $D=0
M2585 877 858 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=145380 $D=0
M2586 878 872 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=136120 $D=0
M2587 879 873 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=140750 $D=0
M2588 880 874 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=145380 $D=0
M2589 163 868 878 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=136120 $D=0
M2590 167 869 879 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=140750 $D=0
M2591 168 870 880 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=145380 $D=0
M2592 883 161 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=136120 $D=0
M2593 884 881 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=140750 $D=0
M2594 885 882 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=145380 $D=0
M2595 881 878 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=136120 $D=0
M2596 882 879 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=140750 $D=0
M2597 162 880 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=145380 $D=0
M2598 163 883 881 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=136120 $D=0
M2599 167 884 882 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=140750 $D=0
M2600 168 885 162 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=145380 $D=0
M2601 888 886 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=136120 $D=0
M2602 889 887 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=140750 $D=0
M2603 890 136 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=145380 $D=0
M2604 163 894 891 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=136120 $D=0
M2605 167 895 892 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=140750 $D=0
M2606 168 896 893 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=145380 $D=0
M2607 897 119 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=136120 $D=0
M2608 898 120 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=140750 $D=0
M2609 899 121 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=145380 $D=0
M2610 894 119 886 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=136120 $D=0
M2611 895 120 887 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=140750 $D=0
M2612 896 121 136 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=145380 $D=0
M2613 888 897 894 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=136120 $D=0
M2614 889 898 895 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=140750 $D=0
M2615 890 899 896 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=145380 $D=0
M2616 900 891 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=136120 $D=0
M2617 901 892 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=140750 $D=0
M2618 902 893 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=145380 $D=0
M2619 164 891 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=136120 $D=0
M2620 886 892 9 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=140750 $D=0
M2621 887 893 136 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=145380 $D=0
M2622 119 900 164 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=136120 $D=0
M2623 120 901 886 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=140750 $D=0
M2624 121 902 887 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=145380 $D=0
M2625 903 164 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=136120 $D=0
M2626 904 886 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=140750 $D=0
M2627 905 887 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=145380 $D=0
M2628 906 891 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=136120 $D=0
M2629 907 892 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=140750 $D=0
M2630 908 893 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=145380 $D=0
M2631 209 891 903 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=136120 $D=0
M2632 210 892 904 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=140750 $D=0
M2633 211 893 905 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=145380 $D=0
M2634 163 906 209 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=136120 $D=0
M2635 9 907 210 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=140750 $D=0
M2636 136 908 211 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=145380 $D=0
M2637 909 165 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=136120 $D=0
M2638 910 165 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=140750 $D=0
M2639 911 165 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=145380 $D=0
M2640 912 165 209 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=136120 $D=0
M2641 913 165 210 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=140750 $D=0
M2642 914 165 211 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=145380 $D=0
M2643 14 909 912 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=136120 $D=0
M2644 15 910 913 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=140750 $D=0
M2645 16 911 914 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=145380 $D=0
M2646 915 166 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=136120 $D=0
M2647 916 166 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=140750 $D=0
M2648 917 166 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=145380 $D=0
M2649 166 166 912 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=136120 $D=0
M2650 166 166 913 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=140750 $D=0
M2651 166 166 914 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=145380 $D=0
M2652 8 915 166 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=136120 $D=0
M2653 9 916 166 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=140750 $D=0
M2654 136 917 166 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=145380 $D=0
M2655 918 114 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=136120 $D=0
M2656 919 114 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=140750 $D=0
M2657 920 114 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=145380 $D=0
M2658 163 918 921 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=136120 $D=0
M2659 167 919 922 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=140750 $D=0
M2660 168 920 923 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=145380 $D=0
M2661 924 114 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=136120 $D=0
M2662 925 114 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=140750 $D=0
M2663 926 114 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=145380 $D=0
M2664 927 921 166 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=136120 $D=0
M2665 928 922 166 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=140750 $D=0
M2666 929 923 166 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=145380 $D=0
M2667 163 927 1071 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=136120 $D=0
M2668 167 928 1072 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=140750 $D=0
M2669 168 929 1073 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=145380 $D=0
M2670 930 1071 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=136120 $D=0
M2671 931 1072 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=140750 $D=0
M2672 932 1073 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=145380 $D=0
M2673 927 918 930 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=136120 $D=0
M2674 928 919 931 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=140750 $D=0
M2675 929 920 932 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=145380 $D=0
M2676 933 924 930 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=136120 $D=0
M2677 934 925 931 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=140750 $D=0
M2678 935 926 932 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=145380 $D=0
M2679 163 939 936 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=136120 $D=0
M2680 167 940 937 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=140750 $D=0
M2681 168 941 938 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=145380 $D=0
M2682 939 114 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=136120 $D=0
M2683 940 114 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=140750 $D=0
M2684 941 114 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=145380 $D=0
M2685 1074 933 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=136120 $D=0
M2686 1075 934 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=140750 $D=0
M2687 1076 935 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=145380 $D=0
M2688 942 939 1074 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=136120 $D=0
M2689 943 940 1075 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=140750 $D=0
M2690 944 941 1076 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=145380 $D=0
M2691 163 942 119 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=136120 $D=0
M2692 167 943 120 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=140750 $D=0
M2693 168 944 121 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=145380 $D=0
M2694 1077 119 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=136120 $D=0
M2695 1078 120 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=140750 $D=0
M2696 1079 121 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=145380 $D=0
M2697 942 936 1077 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=136120 $D=0
M2698 943 937 1078 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=140750 $D=0
M2699 944 938 1079 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=145380 $D=0
.ENDS
***************************************
.SUBCKT ICV_25 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141
+ 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159
** N=787 EP=158 IP=1514 FDC=1800
M0 169 1 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=125610 $D=1
M1 170 1 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=130240 $D=1
M2 171 169 2 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=125610 $D=1
M3 172 170 3 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=130240 $D=1
M4 7 1 171 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=125610 $D=1
M5 8 1 172 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=130240 $D=1
M6 173 169 2 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=125610 $D=1
M7 174 170 3 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=130240 $D=1
M8 2 1 173 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=125610 $D=1
M9 3 1 174 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=130240 $D=1
M10 175 169 2 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=125610 $D=1
M11 176 170 3 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=130240 $D=1
M12 2 1 175 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=125610 $D=1
M13 3 1 176 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=130240 $D=1
M14 179 177 175 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=125610 $D=1
M15 180 178 176 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=130240 $D=1
M16 177 4 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=125610 $D=1
M17 178 4 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=130240 $D=1
M18 181 177 173 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=125610 $D=1
M19 182 178 174 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=130240 $D=1
M20 171 4 181 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=125610 $D=1
M21 172 4 182 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=130240 $D=1
M22 183 5 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=125610 $D=1
M23 184 5 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=130240 $D=1
M24 185 183 181 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=125610 $D=1
M25 186 184 182 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=130240 $D=1
M26 179 5 185 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=125610 $D=1
M27 180 5 186 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=130240 $D=1
M28 187 6 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=125610 $D=1
M29 188 6 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=130240 $D=1
M30 189 187 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=125610 $D=1
M31 190 188 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=130240 $D=1
M32 9 6 189 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=125610 $D=1
M33 10 6 190 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=130240 $D=1
M34 191 187 11 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=125610 $D=1
M35 192 188 12 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=130240 $D=1
M36 193 6 191 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=125610 $D=1
M37 194 6 192 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=130240 $D=1
M38 197 187 195 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=125610 $D=1
M39 198 188 196 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=130240 $D=1
M40 185 6 197 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=125610 $D=1
M41 186 6 198 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=130240 $D=1
M42 201 199 197 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=125610 $D=1
M43 202 200 198 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=130240 $D=1
M44 199 13 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=125610 $D=1
M45 200 13 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=130240 $D=1
M46 203 199 191 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=125610 $D=1
M47 204 200 192 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=130240 $D=1
M48 189 13 203 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=125610 $D=1
M49 190 13 204 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=130240 $D=1
M50 205 14 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=125610 $D=1
M51 206 14 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=130240 $D=1
M52 207 205 203 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=125610 $D=1
M53 208 206 204 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=130240 $D=1
M54 201 14 207 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=125610 $D=1
M55 202 14 208 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=130240 $D=1
M56 7 15 209 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=125610 $D=1
M57 8 15 210 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=130240 $D=1
M58 211 16 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=125610 $D=1
M59 212 16 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=130240 $D=1
M60 213 15 207 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=125610 $D=1
M61 214 15 208 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=130240 $D=1
M62 7 213 680 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=125610 $D=1
M63 8 214 681 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=130240 $D=1
M64 215 680 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=125610 $D=1
M65 216 681 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=130240 $D=1
M66 213 209 215 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=125610 $D=1
M67 214 210 216 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=130240 $D=1
M68 215 16 217 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=125610 $D=1
M69 216 16 218 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=130240 $D=1
M70 221 17 215 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=125610 $D=1
M71 222 17 216 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=130240 $D=1
M72 219 17 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=125610 $D=1
M73 220 17 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=130240 $D=1
M74 7 18 223 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=125610 $D=1
M75 8 18 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=130240 $D=1
M76 225 19 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=125610 $D=1
M77 226 19 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=130240 $D=1
M78 227 18 207 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=125610 $D=1
M79 228 18 208 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=130240 $D=1
M80 7 227 682 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=125610 $D=1
M81 8 228 683 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=130240 $D=1
M82 229 682 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=125610 $D=1
M83 230 683 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=130240 $D=1
M84 227 223 229 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=125610 $D=1
M85 228 224 230 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=130240 $D=1
M86 229 19 217 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=125610 $D=1
M87 230 19 218 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=130240 $D=1
M88 221 20 229 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=125610 $D=1
M89 222 20 230 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=130240 $D=1
M90 231 20 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=125610 $D=1
M91 232 20 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=130240 $D=1
M92 7 21 233 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=125610 $D=1
M93 8 21 234 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=130240 $D=1
M94 235 22 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=125610 $D=1
M95 236 22 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=130240 $D=1
M96 237 21 207 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=125610 $D=1
M97 238 21 208 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=130240 $D=1
M98 7 237 684 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=125610 $D=1
M99 8 238 685 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=130240 $D=1
M100 239 684 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=125610 $D=1
M101 240 685 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=130240 $D=1
M102 237 233 239 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=125610 $D=1
M103 238 234 240 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=130240 $D=1
M104 239 22 217 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=125610 $D=1
M105 240 22 218 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=130240 $D=1
M106 221 23 239 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=125610 $D=1
M107 222 23 240 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=130240 $D=1
M108 241 23 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=125610 $D=1
M109 242 23 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=130240 $D=1
M110 7 24 243 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=125610 $D=1
M111 8 24 244 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=130240 $D=1
M112 245 25 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=125610 $D=1
M113 246 25 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=130240 $D=1
M114 247 24 207 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=125610 $D=1
M115 248 24 208 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=130240 $D=1
M116 7 247 686 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=125610 $D=1
M117 8 248 687 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=130240 $D=1
M118 249 686 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=125610 $D=1
M119 250 687 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=130240 $D=1
M120 247 243 249 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=125610 $D=1
M121 248 244 250 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=130240 $D=1
M122 249 25 217 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=125610 $D=1
M123 250 25 218 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=130240 $D=1
M124 221 26 249 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=125610 $D=1
M125 222 26 250 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=130240 $D=1
M126 251 26 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=125610 $D=1
M127 252 26 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=130240 $D=1
M128 7 27 253 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=125610 $D=1
M129 8 27 254 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=130240 $D=1
M130 255 28 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=125610 $D=1
M131 256 28 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=130240 $D=1
M132 257 27 207 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=125610 $D=1
M133 258 27 208 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=130240 $D=1
M134 7 257 688 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=125610 $D=1
M135 8 258 689 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=130240 $D=1
M136 259 688 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=125610 $D=1
M137 260 689 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=130240 $D=1
M138 257 253 259 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=125610 $D=1
M139 258 254 260 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=130240 $D=1
M140 259 28 217 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=125610 $D=1
M141 260 28 218 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=130240 $D=1
M142 221 29 259 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=125610 $D=1
M143 222 29 260 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=130240 $D=1
M144 261 29 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=125610 $D=1
M145 262 29 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=130240 $D=1
M146 7 30 263 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=125610 $D=1
M147 8 30 264 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=130240 $D=1
M148 265 31 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=125610 $D=1
M149 266 31 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=130240 $D=1
M150 267 30 207 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=125610 $D=1
M151 268 30 208 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=130240 $D=1
M152 7 267 690 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=125610 $D=1
M153 8 268 691 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=130240 $D=1
M154 269 690 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=125610 $D=1
M155 270 691 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=130240 $D=1
M156 267 263 269 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=125610 $D=1
M157 268 264 270 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=130240 $D=1
M158 269 31 217 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=125610 $D=1
M159 270 31 218 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=130240 $D=1
M160 221 32 269 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=125610 $D=1
M161 222 32 270 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=130240 $D=1
M162 271 32 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=125610 $D=1
M163 272 32 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=130240 $D=1
M164 7 33 273 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=125610 $D=1
M165 8 33 274 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=130240 $D=1
M166 275 34 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=125610 $D=1
M167 276 34 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=130240 $D=1
M168 277 33 207 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=125610 $D=1
M169 278 33 208 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=130240 $D=1
M170 7 277 692 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=125610 $D=1
M171 8 278 693 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=130240 $D=1
M172 279 692 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=125610 $D=1
M173 280 693 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=130240 $D=1
M174 277 273 279 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=125610 $D=1
M175 278 274 280 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=130240 $D=1
M176 279 34 217 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=125610 $D=1
M177 280 34 218 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=130240 $D=1
M178 221 35 279 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=125610 $D=1
M179 222 35 280 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=130240 $D=1
M180 281 35 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=125610 $D=1
M181 282 35 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=130240 $D=1
M182 7 36 283 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=125610 $D=1
M183 8 36 284 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=130240 $D=1
M184 285 37 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=125610 $D=1
M185 286 37 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=130240 $D=1
M186 287 36 207 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=125610 $D=1
M187 288 36 208 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=130240 $D=1
M188 7 287 694 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=125610 $D=1
M189 8 288 695 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=130240 $D=1
M190 289 694 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=125610 $D=1
M191 290 695 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=130240 $D=1
M192 287 283 289 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=125610 $D=1
M193 288 284 290 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=130240 $D=1
M194 289 37 217 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=125610 $D=1
M195 290 37 218 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=130240 $D=1
M196 221 38 289 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=125610 $D=1
M197 222 38 290 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=130240 $D=1
M198 291 38 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=125610 $D=1
M199 292 38 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=130240 $D=1
M200 7 39 293 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=125610 $D=1
M201 8 39 294 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=130240 $D=1
M202 295 40 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=125610 $D=1
M203 296 40 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=130240 $D=1
M204 297 39 207 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=125610 $D=1
M205 298 39 208 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=130240 $D=1
M206 7 297 696 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=125610 $D=1
M207 8 298 697 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=130240 $D=1
M208 299 696 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=125610 $D=1
M209 300 697 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=130240 $D=1
M210 297 293 299 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=125610 $D=1
M211 298 294 300 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=130240 $D=1
M212 299 40 217 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=125610 $D=1
M213 300 40 218 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=130240 $D=1
M214 221 41 299 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=125610 $D=1
M215 222 41 300 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=130240 $D=1
M216 301 41 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=125610 $D=1
M217 302 41 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=130240 $D=1
M218 7 42 303 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=125610 $D=1
M219 8 42 304 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=130240 $D=1
M220 305 43 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=125610 $D=1
M221 306 43 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=130240 $D=1
M222 307 42 207 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=125610 $D=1
M223 308 42 208 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=130240 $D=1
M224 7 307 698 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=125610 $D=1
M225 8 308 699 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=130240 $D=1
M226 309 698 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=125610 $D=1
M227 310 699 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=130240 $D=1
M228 307 303 309 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=125610 $D=1
M229 308 304 310 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=130240 $D=1
M230 309 43 217 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=125610 $D=1
M231 310 43 218 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=130240 $D=1
M232 221 44 309 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=125610 $D=1
M233 222 44 310 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=130240 $D=1
M234 311 44 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=125610 $D=1
M235 312 44 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=130240 $D=1
M236 7 45 313 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=125610 $D=1
M237 8 45 314 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=130240 $D=1
M238 315 46 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=125610 $D=1
M239 316 46 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=130240 $D=1
M240 317 45 207 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=125610 $D=1
M241 318 45 208 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=130240 $D=1
M242 7 317 700 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=125610 $D=1
M243 8 318 701 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=130240 $D=1
M244 319 700 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=125610 $D=1
M245 320 701 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=130240 $D=1
M246 317 313 319 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=125610 $D=1
M247 318 314 320 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=130240 $D=1
M248 319 46 217 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=125610 $D=1
M249 320 46 218 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=130240 $D=1
M250 221 47 319 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=125610 $D=1
M251 222 47 320 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=130240 $D=1
M252 321 47 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=125610 $D=1
M253 322 47 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=130240 $D=1
M254 7 48 323 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=125610 $D=1
M255 8 48 324 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=130240 $D=1
M256 325 49 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=125610 $D=1
M257 326 49 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=130240 $D=1
M258 327 48 207 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=125610 $D=1
M259 328 48 208 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=130240 $D=1
M260 7 327 702 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=125610 $D=1
M261 8 328 703 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=130240 $D=1
M262 329 702 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=125610 $D=1
M263 330 703 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=130240 $D=1
M264 327 323 329 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=125610 $D=1
M265 328 324 330 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=130240 $D=1
M266 329 49 217 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=125610 $D=1
M267 330 49 218 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=130240 $D=1
M268 221 50 329 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=125610 $D=1
M269 222 50 330 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=130240 $D=1
M270 331 50 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=125610 $D=1
M271 332 50 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=130240 $D=1
M272 7 51 333 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=125610 $D=1
M273 8 51 334 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=130240 $D=1
M274 335 52 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=125610 $D=1
M275 336 52 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=130240 $D=1
M276 337 51 207 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=125610 $D=1
M277 338 51 208 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=130240 $D=1
M278 7 337 704 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=125610 $D=1
M279 8 338 705 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=130240 $D=1
M280 339 704 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=125610 $D=1
M281 340 705 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=130240 $D=1
M282 337 333 339 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=125610 $D=1
M283 338 334 340 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=130240 $D=1
M284 339 52 217 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=125610 $D=1
M285 340 52 218 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=130240 $D=1
M286 221 53 339 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=125610 $D=1
M287 222 53 340 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=130240 $D=1
M288 341 53 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=125610 $D=1
M289 342 53 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=130240 $D=1
M290 7 54 343 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=125610 $D=1
M291 8 54 344 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=130240 $D=1
M292 345 55 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=125610 $D=1
M293 346 55 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=130240 $D=1
M294 347 54 207 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=125610 $D=1
M295 348 54 208 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=130240 $D=1
M296 7 347 706 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=125610 $D=1
M297 8 348 707 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=130240 $D=1
M298 349 706 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=125610 $D=1
M299 350 707 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=130240 $D=1
M300 347 343 349 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=125610 $D=1
M301 348 344 350 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=130240 $D=1
M302 349 55 217 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=125610 $D=1
M303 350 55 218 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=130240 $D=1
M304 221 56 349 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=125610 $D=1
M305 222 56 350 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=130240 $D=1
M306 351 56 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=125610 $D=1
M307 352 56 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=130240 $D=1
M308 7 57 353 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=125610 $D=1
M309 8 57 354 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=130240 $D=1
M310 355 58 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=125610 $D=1
M311 356 58 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=130240 $D=1
M312 357 57 207 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=125610 $D=1
M313 358 57 208 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=130240 $D=1
M314 7 357 708 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=125610 $D=1
M315 8 358 709 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=130240 $D=1
M316 359 708 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=125610 $D=1
M317 360 709 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=130240 $D=1
M318 357 353 359 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=125610 $D=1
M319 358 354 360 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=130240 $D=1
M320 359 58 217 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=125610 $D=1
M321 360 58 218 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=130240 $D=1
M322 221 59 359 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=125610 $D=1
M323 222 59 360 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=130240 $D=1
M324 361 59 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=125610 $D=1
M325 362 59 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=130240 $D=1
M326 7 60 363 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=125610 $D=1
M327 8 60 364 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=130240 $D=1
M328 365 61 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=125610 $D=1
M329 366 61 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=130240 $D=1
M330 367 60 207 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=125610 $D=1
M331 368 60 208 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=130240 $D=1
M332 7 367 710 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=125610 $D=1
M333 8 368 711 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=130240 $D=1
M334 369 710 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=125610 $D=1
M335 370 711 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=130240 $D=1
M336 367 363 369 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=125610 $D=1
M337 368 364 370 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=130240 $D=1
M338 369 61 217 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=125610 $D=1
M339 370 61 218 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=130240 $D=1
M340 221 62 369 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=125610 $D=1
M341 222 62 370 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=130240 $D=1
M342 371 62 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=125610 $D=1
M343 372 62 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=130240 $D=1
M344 7 63 373 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=125610 $D=1
M345 8 63 374 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=130240 $D=1
M346 375 64 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=125610 $D=1
M347 376 64 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=130240 $D=1
M348 377 63 207 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=125610 $D=1
M349 378 63 208 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=130240 $D=1
M350 7 377 712 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=125610 $D=1
M351 8 378 713 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=130240 $D=1
M352 379 712 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=125610 $D=1
M353 380 713 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=130240 $D=1
M354 377 373 379 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=125610 $D=1
M355 378 374 380 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=130240 $D=1
M356 379 64 217 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=125610 $D=1
M357 380 64 218 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=130240 $D=1
M358 221 65 379 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=125610 $D=1
M359 222 65 380 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=130240 $D=1
M360 381 65 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=125610 $D=1
M361 382 65 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=130240 $D=1
M362 7 66 383 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=125610 $D=1
M363 8 66 384 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=130240 $D=1
M364 385 67 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=125610 $D=1
M365 386 67 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=130240 $D=1
M366 387 66 207 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=125610 $D=1
M367 388 66 208 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=130240 $D=1
M368 7 387 714 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=125610 $D=1
M369 8 388 715 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=130240 $D=1
M370 389 714 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=125610 $D=1
M371 390 715 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=130240 $D=1
M372 387 383 389 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=125610 $D=1
M373 388 384 390 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=130240 $D=1
M374 389 67 217 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=125610 $D=1
M375 390 67 218 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=130240 $D=1
M376 221 68 389 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=125610 $D=1
M377 222 68 390 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=130240 $D=1
M378 391 68 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=125610 $D=1
M379 392 68 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=130240 $D=1
M380 7 69 393 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=125610 $D=1
M381 8 69 394 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=130240 $D=1
M382 395 70 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=125610 $D=1
M383 396 70 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=130240 $D=1
M384 397 69 207 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=125610 $D=1
M385 398 69 208 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=130240 $D=1
M386 7 397 716 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=125610 $D=1
M387 8 398 717 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=130240 $D=1
M388 399 716 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=125610 $D=1
M389 400 717 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=130240 $D=1
M390 397 393 399 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=125610 $D=1
M391 398 394 400 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=130240 $D=1
M392 399 70 217 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=125610 $D=1
M393 400 70 218 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=130240 $D=1
M394 221 71 399 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=125610 $D=1
M395 222 71 400 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=130240 $D=1
M396 401 71 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=125610 $D=1
M397 402 71 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=130240 $D=1
M398 7 72 403 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=125610 $D=1
M399 8 72 404 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=130240 $D=1
M400 405 73 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=125610 $D=1
M401 406 73 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=130240 $D=1
M402 407 72 207 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=125610 $D=1
M403 408 72 208 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=130240 $D=1
M404 7 407 718 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=125610 $D=1
M405 8 408 719 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=130240 $D=1
M406 409 718 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=125610 $D=1
M407 410 719 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=130240 $D=1
M408 407 403 409 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=125610 $D=1
M409 408 404 410 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=130240 $D=1
M410 409 73 217 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=125610 $D=1
M411 410 73 218 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=130240 $D=1
M412 221 74 409 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=125610 $D=1
M413 222 74 410 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=130240 $D=1
M414 411 74 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=125610 $D=1
M415 412 74 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=130240 $D=1
M416 7 75 413 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=125610 $D=1
M417 8 75 414 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=130240 $D=1
M418 415 76 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=125610 $D=1
M419 416 76 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=130240 $D=1
M420 417 75 207 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=125610 $D=1
M421 418 75 208 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=130240 $D=1
M422 7 417 720 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=125610 $D=1
M423 8 418 721 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=130240 $D=1
M424 419 720 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=125610 $D=1
M425 420 721 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=130240 $D=1
M426 417 413 419 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=125610 $D=1
M427 418 414 420 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=130240 $D=1
M428 419 76 217 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=125610 $D=1
M429 420 76 218 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=130240 $D=1
M430 221 77 419 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=125610 $D=1
M431 222 77 420 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=130240 $D=1
M432 421 77 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=125610 $D=1
M433 422 77 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=130240 $D=1
M434 7 78 423 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=125610 $D=1
M435 8 78 424 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=130240 $D=1
M436 425 79 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=125610 $D=1
M437 426 79 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=130240 $D=1
M438 427 78 207 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=125610 $D=1
M439 428 78 208 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=130240 $D=1
M440 7 427 722 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=125610 $D=1
M441 8 428 723 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=130240 $D=1
M442 429 722 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=125610 $D=1
M443 430 723 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=130240 $D=1
M444 427 423 429 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=125610 $D=1
M445 428 424 430 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=130240 $D=1
M446 429 79 217 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=125610 $D=1
M447 430 79 218 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=130240 $D=1
M448 221 80 429 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=125610 $D=1
M449 222 80 430 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=130240 $D=1
M450 431 80 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=125610 $D=1
M451 432 80 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=130240 $D=1
M452 7 81 433 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=125610 $D=1
M453 8 81 434 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=130240 $D=1
M454 435 82 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=125610 $D=1
M455 436 82 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=130240 $D=1
M456 437 81 207 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=125610 $D=1
M457 438 81 208 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=130240 $D=1
M458 7 437 724 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=125610 $D=1
M459 8 438 725 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=130240 $D=1
M460 439 724 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=125610 $D=1
M461 440 725 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=130240 $D=1
M462 437 433 439 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=125610 $D=1
M463 438 434 440 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=130240 $D=1
M464 439 82 217 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=125610 $D=1
M465 440 82 218 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=130240 $D=1
M466 221 83 439 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=125610 $D=1
M467 222 83 440 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=130240 $D=1
M468 441 83 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=125610 $D=1
M469 442 83 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=130240 $D=1
M470 7 84 443 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=125610 $D=1
M471 8 84 444 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=130240 $D=1
M472 445 85 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=125610 $D=1
M473 446 85 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=130240 $D=1
M474 447 84 207 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=125610 $D=1
M475 448 84 208 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=130240 $D=1
M476 7 447 726 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=125610 $D=1
M477 8 448 727 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=130240 $D=1
M478 449 726 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=125610 $D=1
M479 450 727 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=130240 $D=1
M480 447 443 449 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=125610 $D=1
M481 448 444 450 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=130240 $D=1
M482 449 85 217 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=125610 $D=1
M483 450 85 218 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=130240 $D=1
M484 221 86 449 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=125610 $D=1
M485 222 86 450 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=130240 $D=1
M486 451 86 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=125610 $D=1
M487 452 86 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=130240 $D=1
M488 7 87 453 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=125610 $D=1
M489 8 87 454 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=130240 $D=1
M490 455 88 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=125610 $D=1
M491 456 88 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=130240 $D=1
M492 457 87 207 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=125610 $D=1
M493 458 87 208 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=130240 $D=1
M494 7 457 728 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=125610 $D=1
M495 8 458 729 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=130240 $D=1
M496 459 728 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=125610 $D=1
M497 460 729 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=130240 $D=1
M498 457 453 459 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=125610 $D=1
M499 458 454 460 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=130240 $D=1
M500 459 88 217 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=125610 $D=1
M501 460 88 218 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=130240 $D=1
M502 221 89 459 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=125610 $D=1
M503 222 89 460 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=130240 $D=1
M504 461 89 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=125610 $D=1
M505 462 89 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=130240 $D=1
M506 7 90 463 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=125610 $D=1
M507 8 90 464 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=130240 $D=1
M508 465 91 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=125610 $D=1
M509 466 91 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=130240 $D=1
M510 467 90 207 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=125610 $D=1
M511 468 90 208 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=130240 $D=1
M512 7 467 730 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=125610 $D=1
M513 8 468 731 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=130240 $D=1
M514 469 730 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=125610 $D=1
M515 470 731 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=130240 $D=1
M516 467 463 469 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=125610 $D=1
M517 468 464 470 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=130240 $D=1
M518 469 91 217 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=125610 $D=1
M519 470 91 218 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=130240 $D=1
M520 221 92 469 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=125610 $D=1
M521 222 92 470 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=130240 $D=1
M522 471 92 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=125610 $D=1
M523 472 92 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=130240 $D=1
M524 7 93 473 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=125610 $D=1
M525 8 93 474 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=130240 $D=1
M526 475 94 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=125610 $D=1
M527 476 94 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=130240 $D=1
M528 477 93 207 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=125610 $D=1
M529 478 93 208 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=130240 $D=1
M530 7 477 732 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=125610 $D=1
M531 8 478 733 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=130240 $D=1
M532 479 732 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=125610 $D=1
M533 480 733 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=130240 $D=1
M534 477 473 479 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=125610 $D=1
M535 478 474 480 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=130240 $D=1
M536 479 94 217 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=125610 $D=1
M537 480 94 218 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=130240 $D=1
M538 221 95 479 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=125610 $D=1
M539 222 95 480 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=130240 $D=1
M540 481 95 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=125610 $D=1
M541 482 95 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=130240 $D=1
M542 7 96 483 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=125610 $D=1
M543 8 96 484 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=130240 $D=1
M544 485 97 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=125610 $D=1
M545 486 97 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=130240 $D=1
M546 487 96 207 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=125610 $D=1
M547 488 96 208 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=130240 $D=1
M548 7 487 734 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=125610 $D=1
M549 8 488 735 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=130240 $D=1
M550 489 734 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=125610 $D=1
M551 490 735 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=130240 $D=1
M552 487 483 489 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=125610 $D=1
M553 488 484 490 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=130240 $D=1
M554 489 97 217 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=125610 $D=1
M555 490 97 218 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=130240 $D=1
M556 221 98 489 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=125610 $D=1
M557 222 98 490 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=130240 $D=1
M558 491 98 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=125610 $D=1
M559 492 98 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=130240 $D=1
M560 7 99 493 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=125610 $D=1
M561 8 99 494 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=130240 $D=1
M562 495 100 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=125610 $D=1
M563 496 100 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=130240 $D=1
M564 497 99 207 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=125610 $D=1
M565 498 99 208 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=130240 $D=1
M566 7 497 736 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=125610 $D=1
M567 8 498 737 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=130240 $D=1
M568 499 736 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=125610 $D=1
M569 500 737 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=130240 $D=1
M570 497 493 499 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=125610 $D=1
M571 498 494 500 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=130240 $D=1
M572 499 100 217 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=125610 $D=1
M573 500 100 218 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=130240 $D=1
M574 221 101 499 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=125610 $D=1
M575 222 101 500 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=130240 $D=1
M576 501 101 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=125610 $D=1
M577 502 101 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=130240 $D=1
M578 7 102 503 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=125610 $D=1
M579 8 102 504 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=130240 $D=1
M580 505 103 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=125610 $D=1
M581 506 103 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=130240 $D=1
M582 507 102 207 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=125610 $D=1
M583 508 102 208 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=130240 $D=1
M584 7 507 738 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=125610 $D=1
M585 8 508 739 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=130240 $D=1
M586 509 738 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=125610 $D=1
M587 510 739 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=130240 $D=1
M588 507 503 509 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=125610 $D=1
M589 508 504 510 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=130240 $D=1
M590 509 103 217 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=125610 $D=1
M591 510 103 218 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=130240 $D=1
M592 221 104 509 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=125610 $D=1
M593 222 104 510 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=130240 $D=1
M594 511 104 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=125610 $D=1
M595 512 104 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=130240 $D=1
M596 7 105 513 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=125610 $D=1
M597 8 105 514 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=130240 $D=1
M598 515 106 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=125610 $D=1
M599 516 106 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=130240 $D=1
M600 517 105 207 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=125610 $D=1
M601 518 105 208 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=130240 $D=1
M602 7 517 740 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=125610 $D=1
M603 8 518 741 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=130240 $D=1
M604 519 740 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=125610 $D=1
M605 520 741 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=130240 $D=1
M606 517 513 519 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=125610 $D=1
M607 518 514 520 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=130240 $D=1
M608 519 106 217 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=125610 $D=1
M609 520 106 218 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=130240 $D=1
M610 221 107 519 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=125610 $D=1
M611 222 107 520 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=130240 $D=1
M612 521 107 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=125610 $D=1
M613 522 107 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=130240 $D=1
M614 7 108 523 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=125610 $D=1
M615 8 108 524 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=130240 $D=1
M616 525 109 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=125610 $D=1
M617 526 109 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=130240 $D=1
M618 7 109 217 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=125610 $D=1
M619 8 109 218 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=130240 $D=1
M620 221 108 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=125610 $D=1
M621 222 108 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=130240 $D=1
M622 7 529 527 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=125610 $D=1
M623 8 530 528 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=130240 $D=1
M624 529 110 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=125610 $D=1
M625 530 110 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=130240 $D=1
M626 742 217 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=125610 $D=1
M627 743 218 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=130240 $D=1
M628 531 527 742 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=125610 $D=1
M629 532 528 743 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=130240 $D=1
M630 7 531 533 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=125610 $D=1
M631 8 532 534 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=130240 $D=1
M632 744 533 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=125610 $D=1
M633 745 534 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=130240 $D=1
M634 531 529 744 7 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=125610 $D=1
M635 532 530 745 8 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=130240 $D=1
M636 7 537 535 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=125610 $D=1
M637 8 538 536 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=130240 $D=1
M638 537 110 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=125610 $D=1
M639 538 110 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=130240 $D=1
M640 746 221 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=125610 $D=1
M641 747 222 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=130240 $D=1
M642 539 535 746 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=125610 $D=1
M643 540 536 747 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=130240 $D=1
M644 7 539 111 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=125610 $D=1
M645 8 540 112 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=130240 $D=1
M646 748 111 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=125610 $D=1
M647 749 112 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=130240 $D=1
M648 539 537 748 7 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=125610 $D=1
M649 540 538 749 8 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=130240 $D=1
M650 541 113 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=125610 $D=1
M651 542 113 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=130240 $D=1
M652 543 541 533 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=125610 $D=1
M653 544 542 534 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=130240 $D=1
M654 114 113 543 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=125610 $D=1
M655 115 113 544 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=130240 $D=1
M656 545 116 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=125610 $D=1
M657 546 116 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=130240 $D=1
M658 547 545 111 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=125610 $D=1
M659 548 546 112 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=130240 $D=1
M660 750 116 547 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=125610 $D=1
M661 751 116 548 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=130240 $D=1
M662 7 111 750 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=125610 $D=1
M663 8 112 751 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=130240 $D=1
M664 549 117 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=125610 $D=1
M665 550 117 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=130240 $D=1
M666 118 549 547 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=125610 $D=1
M667 119 550 548 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=130240 $D=1
M668 9 117 118 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=125610 $D=1
M669 10 117 119 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=130240 $D=1
M670 552 551 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=125610 $D=1
M671 553 120 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=130240 $D=1
M672 7 556 554 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=125610 $D=1
M673 8 557 555 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=130240 $D=1
M674 558 543 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=125610 $D=1
M675 559 544 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=130240 $D=1
M676 556 558 551 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=125610 $D=1
M677 557 559 120 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=130240 $D=1
M678 552 543 556 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=125610 $D=1
M679 553 544 557 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=130240 $D=1
M680 560 554 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=125610 $D=1
M681 561 555 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=130240 $D=1
M682 562 560 118 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=125610 $D=1
M683 551 561 119 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=130240 $D=1
M684 543 554 562 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=125610 $D=1
M685 544 555 551 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=130240 $D=1
M686 563 562 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=125610 $D=1
M687 564 551 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=130240 $D=1
M688 565 554 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=125610 $D=1
M689 566 555 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=130240 $D=1
M690 567 565 563 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=125610 $D=1
M691 568 566 564 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=130240 $D=1
M692 118 554 567 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=125610 $D=1
M693 119 555 568 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=130240 $D=1
M694 569 543 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=125610 $D=1
M695 570 544 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=130240 $D=1
M696 7 118 569 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=125610 $D=1
M697 8 119 570 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=130240 $D=1
M698 571 567 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=125610 $D=1
M699 572 568 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=130240 $D=1
M700 776 543 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=125610 $D=1
M701 777 544 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=130240 $D=1
M702 573 118 776 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=125610 $D=1
M703 574 119 777 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=130240 $D=1
M704 778 543 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=125610 $D=1
M705 779 544 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=130240 $D=1
M706 575 118 778 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=125610 $D=1
M707 576 119 779 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=130240 $D=1
M708 579 543 577 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=125610 $D=1
M709 580 544 578 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=130240 $D=1
M710 577 118 579 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=125610 $D=1
M711 578 119 580 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=130240 $D=1
M712 7 575 577 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=125610 $D=1
M713 8 576 578 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=130240 $D=1
M714 581 124 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=125610 $D=1
M715 582 124 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=130240 $D=1
M716 583 581 569 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=125610 $D=1
M717 584 582 570 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=130240 $D=1
M718 573 124 583 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=125610 $D=1
M719 574 124 584 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=130240 $D=1
M720 585 581 571 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=125610 $D=1
M721 586 582 572 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=130240 $D=1
M722 579 124 585 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=125610 $D=1
M723 580 124 586 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=130240 $D=1
M724 587 125 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=125610 $D=1
M725 588 125 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=130240 $D=1
M726 589 587 585 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=125610 $D=1
M727 590 588 586 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=130240 $D=1
M728 583 125 589 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=125610 $D=1
M729 584 125 590 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=130240 $D=1
M730 11 589 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=125610 $D=1
M731 12 590 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=130240 $D=1
M732 591 127 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=125610 $D=1
M733 592 127 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=130240 $D=1
M734 593 591 128 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=125610 $D=1
M735 594 592 129 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=130240 $D=1
M736 130 127 593 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=125610 $D=1
M737 118 127 594 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=130240 $D=1
M738 595 127 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=125610 $D=1
M739 596 127 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=130240 $D=1
M740 598 595 131 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=125610 $D=1
M741 599 596 133 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=130240 $D=1
M742 134 127 598 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=125610 $D=1
M743 132 127 599 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=130240 $D=1
M744 600 127 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=125610 $D=1
M745 601 127 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=130240 $D=1
M746 135 600 121 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=125610 $D=1
M747 135 601 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=130240 $D=1
M748 126 127 135 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=125610 $D=1
M749 136 127 135 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=130240 $D=1
M750 602 127 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=125610 $D=1
M751 603 127 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=130240 $D=1
M752 604 602 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=125610 $D=1
M753 605 603 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=130240 $D=1
M754 137 127 604 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=125610 $D=1
M755 138 127 605 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=130240 $D=1
M756 606 127 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=125610 $D=1
M757 607 127 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=130240 $D=1
M758 608 606 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=125610 $D=1
M759 609 607 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=130240 $D=1
M760 139 127 608 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=125610 $D=1
M761 140 127 609 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=130240 $D=1
M762 7 543 758 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=125610 $D=1
M763 8 544 759 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=130240 $D=1
M764 118 758 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=125610 $D=1
M765 128 759 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=130240 $D=1
M766 610 141 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=125610 $D=1
M767 611 141 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=130240 $D=1
M768 142 610 118 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=125610 $D=1
M769 143 611 128 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=130240 $D=1
M770 593 141 142 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=125610 $D=1
M771 594 141 143 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=130240 $D=1
M772 612 144 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=125610 $D=1
M773 613 144 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=130240 $D=1
M774 145 612 142 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=125610 $D=1
M775 123 613 143 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=130240 $D=1
M776 598 144 145 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=125610 $D=1
M777 599 144 123 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=130240 $D=1
M778 614 129 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=125610 $D=1
M779 615 129 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=130240 $D=1
M780 146 614 145 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=125610 $D=1
M781 147 615 123 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=130240 $D=1
M782 135 129 146 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=125610 $D=1
M783 135 129 147 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=130240 $D=1
M784 616 119 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=125610 $D=1
M785 617 119 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=130240 $D=1
M786 148 616 146 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=125610 $D=1
M787 149 617 147 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=130240 $D=1
M788 604 119 148 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=125610 $D=1
M789 605 119 149 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=130240 $D=1
M790 618 118 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=125610 $D=1
M791 619 118 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=130240 $D=1
M792 193 618 148 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=125610 $D=1
M793 194 619 149 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=130240 $D=1
M794 608 118 193 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=125610 $D=1
M795 609 118 194 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=130240 $D=1
M796 620 150 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=125610 $D=1
M797 621 150 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=130240 $D=1
M798 622 620 111 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=125610 $D=1
M799 623 621 112 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=130240 $D=1
M800 9 150 622 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=125610 $D=1
M801 10 150 623 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=130240 $D=1
M802 780 533 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=125610 $D=1
M803 781 534 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=130240 $D=1
M804 624 622 780 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=125610 $D=1
M805 625 623 781 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=130240 $D=1
M806 628 533 626 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=125610 $D=1
M807 629 534 627 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=130240 $D=1
M808 626 622 628 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=125610 $D=1
M809 627 623 629 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=130240 $D=1
M810 7 624 626 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=125610 $D=1
M811 8 625 627 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=130240 $D=1
M812 782 630 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=125610 $D=1
M813 783 631 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=130240 $D=1
M814 760 628 782 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=125610 $D=1
M815 761 629 783 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=130240 $D=1
M816 631 760 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=125610 $D=1
M817 151 761 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=130240 $D=1
M818 632 533 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=125610 $D=1
M819 633 534 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=130240 $D=1
M820 7 634 632 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=125610 $D=1
M821 8 635 633 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=130240 $D=1
M822 634 622 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=125610 $D=1
M823 635 623 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=130240 $D=1
M824 784 632 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=125610 $D=1
M825 785 633 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=130240 $D=1
M826 636 630 784 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=125610 $D=1
M827 637 631 785 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=130240 $D=1
M828 639 152 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=125610 $D=1
M829 640 638 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=130240 $D=1
M830 786 636 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=125610 $D=1
M831 787 637 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=130240 $D=1
M832 638 639 786 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=125610 $D=1
M833 153 640 787 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=130240 $D=1
M834 642 641 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=125610 $D=1
M835 643 154 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=130240 $D=1
M836 7 646 644 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=125610 $D=1
M837 8 647 645 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=130240 $D=1
M838 648 114 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=125610 $D=1
M839 649 115 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=130240 $D=1
M840 646 648 641 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=125610 $D=1
M841 647 649 154 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=130240 $D=1
M842 642 114 646 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=125610 $D=1
M843 643 115 647 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=130240 $D=1
M844 650 644 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=125610 $D=1
M845 651 645 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=130240 $D=1
M846 155 650 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=125610 $D=1
M847 641 651 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=130240 $D=1
M848 114 644 155 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=125610 $D=1
M849 115 645 641 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=130240 $D=1
M850 652 155 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=125610 $D=1
M851 653 641 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=130240 $D=1
M852 654 644 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=125610 $D=1
M853 655 645 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=130240 $D=1
M854 195 654 652 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=125610 $D=1
M855 196 655 653 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=130240 $D=1
M856 7 644 195 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=125610 $D=1
M857 8 645 196 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=130240 $D=1
M858 656 156 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=125610 $D=1
M859 657 156 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=130240 $D=1
M860 658 656 195 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=125610 $D=1
M861 659 657 196 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=130240 $D=1
M862 11 156 658 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=125610 $D=1
M863 12 156 659 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=130240 $D=1
M864 660 157 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=125610 $D=1
M865 661 157 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=130240 $D=1
M866 157 660 658 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=125610 $D=1
M867 157 661 659 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=130240 $D=1
M868 7 157 157 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=125610 $D=1
M869 8 157 157 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=130240 $D=1
M870 662 110 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=125610 $D=1
M871 663 110 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=130240 $D=1
M872 7 662 664 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=125610 $D=1
M873 8 663 665 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=130240 $D=1
M874 666 110 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=125610 $D=1
M875 667 110 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=130240 $D=1
M876 668 662 157 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=125610 $D=1
M877 669 663 157 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=130240 $D=1
M878 7 668 762 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=125610 $D=1
M879 8 669 763 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=130240 $D=1
M880 670 762 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=125610 $D=1
M881 671 763 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=130240 $D=1
M882 668 664 670 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=125610 $D=1
M883 669 665 671 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=130240 $D=1
M884 672 110 670 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=125610 $D=1
M885 673 110 671 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=130240 $D=1
M886 7 676 674 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=125610 $D=1
M887 8 677 675 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=130240 $D=1
M888 676 110 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=125610 $D=1
M889 677 110 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=130240 $D=1
M890 764 672 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=125610 $D=1
M891 765 673 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=130240 $D=1
M892 678 674 764 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=125610 $D=1
M893 679 675 765 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=130240 $D=1
M894 7 678 114 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=125610 $D=1
M895 8 679 115 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=130240 $D=1
M896 766 114 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=125610 $D=1
M897 767 115 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=130240 $D=1
M898 678 676 766 7 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=125610 $D=1
M899 679 677 767 8 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=130240 $D=1
M900 169 1 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=126860 $D=0
M901 170 1 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=131490 $D=0
M902 171 1 2 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=126860 $D=0
M903 172 1 3 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=131490 $D=0
M904 7 169 171 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=126860 $D=0
M905 8 170 172 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=131490 $D=0
M906 173 1 2 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=126860 $D=0
M907 174 1 3 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=131490 $D=0
M908 2 169 173 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=126860 $D=0
M909 3 170 174 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=131490 $D=0
M910 175 1 2 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=126860 $D=0
M911 176 1 3 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=131490 $D=0
M912 2 169 175 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=126860 $D=0
M913 3 170 176 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=131490 $D=0
M914 179 4 175 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=126860 $D=0
M915 180 4 176 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=131490 $D=0
M916 177 4 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=126860 $D=0
M917 178 4 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=131490 $D=0
M918 181 4 173 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=126860 $D=0
M919 182 4 174 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=131490 $D=0
M920 171 177 181 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=126860 $D=0
M921 172 178 182 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=131490 $D=0
M922 183 5 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=126860 $D=0
M923 184 5 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=131490 $D=0
M924 185 5 181 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=126860 $D=0
M925 186 5 182 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=131490 $D=0
M926 179 183 185 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=126860 $D=0
M927 180 184 186 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=131490 $D=0
M928 187 6 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=126860 $D=0
M929 188 6 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=131490 $D=0
M930 189 6 7 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=126860 $D=0
M931 190 6 8 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=131490 $D=0
M932 9 187 189 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=126860 $D=0
M933 10 188 190 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=131490 $D=0
M934 191 6 11 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=126860 $D=0
M935 192 6 12 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=131490 $D=0
M936 193 187 191 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=126860 $D=0
M937 194 188 192 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=131490 $D=0
M938 197 6 195 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=126860 $D=0
M939 198 6 196 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=131490 $D=0
M940 185 187 197 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=126860 $D=0
M941 186 188 198 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=131490 $D=0
M942 201 13 197 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=126860 $D=0
M943 202 13 198 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=131490 $D=0
M944 199 13 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=126860 $D=0
M945 200 13 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=131490 $D=0
M946 203 13 191 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=126860 $D=0
M947 204 13 192 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=131490 $D=0
M948 189 199 203 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=126860 $D=0
M949 190 200 204 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=131490 $D=0
M950 205 14 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=126860 $D=0
M951 206 14 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=131490 $D=0
M952 207 14 203 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=126860 $D=0
M953 208 14 204 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=131490 $D=0
M954 201 205 207 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=126860 $D=0
M955 202 206 208 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=131490 $D=0
M956 158 15 209 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=126860 $D=0
M957 159 15 210 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=131490 $D=0
M958 211 16 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=126860 $D=0
M959 212 16 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=131490 $D=0
M960 213 209 207 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=126860 $D=0
M961 214 210 208 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=131490 $D=0
M962 158 213 680 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=126860 $D=0
M963 159 214 681 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=131490 $D=0
M964 215 680 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=126860 $D=0
M965 216 681 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=131490 $D=0
M966 213 15 215 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=126860 $D=0
M967 214 15 216 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=131490 $D=0
M968 215 211 217 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=126860 $D=0
M969 216 212 218 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=131490 $D=0
M970 221 219 215 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=126860 $D=0
M971 222 220 216 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=131490 $D=0
M972 219 17 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=126860 $D=0
M973 220 17 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=131490 $D=0
M974 158 18 223 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=126860 $D=0
M975 159 18 224 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=131490 $D=0
M976 225 19 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=126860 $D=0
M977 226 19 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=131490 $D=0
M978 227 223 207 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=126860 $D=0
M979 228 224 208 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=131490 $D=0
M980 158 227 682 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=126860 $D=0
M981 159 228 683 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=131490 $D=0
M982 229 682 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=126860 $D=0
M983 230 683 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=131490 $D=0
M984 227 18 229 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=126860 $D=0
M985 228 18 230 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=131490 $D=0
M986 229 225 217 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=126860 $D=0
M987 230 226 218 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=131490 $D=0
M988 221 231 229 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=126860 $D=0
M989 222 232 230 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=131490 $D=0
M990 231 20 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=126860 $D=0
M991 232 20 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=131490 $D=0
M992 158 21 233 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=126860 $D=0
M993 159 21 234 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=131490 $D=0
M994 235 22 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=126860 $D=0
M995 236 22 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=131490 $D=0
M996 237 233 207 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=126860 $D=0
M997 238 234 208 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=131490 $D=0
M998 158 237 684 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=126860 $D=0
M999 159 238 685 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=131490 $D=0
M1000 239 684 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=126860 $D=0
M1001 240 685 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=131490 $D=0
M1002 237 21 239 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=126860 $D=0
M1003 238 21 240 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=131490 $D=0
M1004 239 235 217 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=126860 $D=0
M1005 240 236 218 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=131490 $D=0
M1006 221 241 239 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=126860 $D=0
M1007 222 242 240 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=131490 $D=0
M1008 241 23 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=126860 $D=0
M1009 242 23 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=131490 $D=0
M1010 158 24 243 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=126860 $D=0
M1011 159 24 244 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=131490 $D=0
M1012 245 25 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=126860 $D=0
M1013 246 25 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=131490 $D=0
M1014 247 243 207 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=126860 $D=0
M1015 248 244 208 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=131490 $D=0
M1016 158 247 686 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=126860 $D=0
M1017 159 248 687 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=131490 $D=0
M1018 249 686 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=126860 $D=0
M1019 250 687 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=131490 $D=0
M1020 247 24 249 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=126860 $D=0
M1021 248 24 250 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=131490 $D=0
M1022 249 245 217 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=126860 $D=0
M1023 250 246 218 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=131490 $D=0
M1024 221 251 249 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=126860 $D=0
M1025 222 252 250 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=131490 $D=0
M1026 251 26 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=126860 $D=0
M1027 252 26 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=131490 $D=0
M1028 158 27 253 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=126860 $D=0
M1029 159 27 254 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=131490 $D=0
M1030 255 28 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=126860 $D=0
M1031 256 28 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=131490 $D=0
M1032 257 253 207 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=126860 $D=0
M1033 258 254 208 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=131490 $D=0
M1034 158 257 688 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=126860 $D=0
M1035 159 258 689 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=131490 $D=0
M1036 259 688 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=126860 $D=0
M1037 260 689 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=131490 $D=0
M1038 257 27 259 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=126860 $D=0
M1039 258 27 260 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=131490 $D=0
M1040 259 255 217 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=126860 $D=0
M1041 260 256 218 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=131490 $D=0
M1042 221 261 259 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=126860 $D=0
M1043 222 262 260 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=131490 $D=0
M1044 261 29 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=126860 $D=0
M1045 262 29 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=131490 $D=0
M1046 158 30 263 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=126860 $D=0
M1047 159 30 264 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=131490 $D=0
M1048 265 31 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=126860 $D=0
M1049 266 31 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=131490 $D=0
M1050 267 263 207 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=126860 $D=0
M1051 268 264 208 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=131490 $D=0
M1052 158 267 690 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=126860 $D=0
M1053 159 268 691 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=131490 $D=0
M1054 269 690 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=126860 $D=0
M1055 270 691 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=131490 $D=0
M1056 267 30 269 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=126860 $D=0
M1057 268 30 270 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=131490 $D=0
M1058 269 265 217 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=126860 $D=0
M1059 270 266 218 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=131490 $D=0
M1060 221 271 269 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=126860 $D=0
M1061 222 272 270 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=131490 $D=0
M1062 271 32 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=126860 $D=0
M1063 272 32 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=131490 $D=0
M1064 158 33 273 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=126860 $D=0
M1065 159 33 274 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=131490 $D=0
M1066 275 34 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=126860 $D=0
M1067 276 34 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=131490 $D=0
M1068 277 273 207 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=126860 $D=0
M1069 278 274 208 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=131490 $D=0
M1070 158 277 692 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=126860 $D=0
M1071 159 278 693 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=131490 $D=0
M1072 279 692 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=126860 $D=0
M1073 280 693 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=131490 $D=0
M1074 277 33 279 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=126860 $D=0
M1075 278 33 280 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=131490 $D=0
M1076 279 275 217 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=126860 $D=0
M1077 280 276 218 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=131490 $D=0
M1078 221 281 279 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=126860 $D=0
M1079 222 282 280 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=131490 $D=0
M1080 281 35 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=126860 $D=0
M1081 282 35 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=131490 $D=0
M1082 158 36 283 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=126860 $D=0
M1083 159 36 284 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=131490 $D=0
M1084 285 37 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=126860 $D=0
M1085 286 37 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=131490 $D=0
M1086 287 283 207 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=126860 $D=0
M1087 288 284 208 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=131490 $D=0
M1088 158 287 694 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=126860 $D=0
M1089 159 288 695 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=131490 $D=0
M1090 289 694 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=126860 $D=0
M1091 290 695 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=131490 $D=0
M1092 287 36 289 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=126860 $D=0
M1093 288 36 290 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=131490 $D=0
M1094 289 285 217 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=126860 $D=0
M1095 290 286 218 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=131490 $D=0
M1096 221 291 289 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=126860 $D=0
M1097 222 292 290 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=131490 $D=0
M1098 291 38 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=126860 $D=0
M1099 292 38 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=131490 $D=0
M1100 158 39 293 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=126860 $D=0
M1101 159 39 294 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=131490 $D=0
M1102 295 40 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=126860 $D=0
M1103 296 40 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=131490 $D=0
M1104 297 293 207 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=126860 $D=0
M1105 298 294 208 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=131490 $D=0
M1106 158 297 696 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=126860 $D=0
M1107 159 298 697 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=131490 $D=0
M1108 299 696 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=126860 $D=0
M1109 300 697 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=131490 $D=0
M1110 297 39 299 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=126860 $D=0
M1111 298 39 300 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=131490 $D=0
M1112 299 295 217 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=126860 $D=0
M1113 300 296 218 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=131490 $D=0
M1114 221 301 299 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=126860 $D=0
M1115 222 302 300 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=131490 $D=0
M1116 301 41 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=126860 $D=0
M1117 302 41 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=131490 $D=0
M1118 158 42 303 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=126860 $D=0
M1119 159 42 304 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=131490 $D=0
M1120 305 43 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=126860 $D=0
M1121 306 43 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=131490 $D=0
M1122 307 303 207 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=126860 $D=0
M1123 308 304 208 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=131490 $D=0
M1124 158 307 698 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=126860 $D=0
M1125 159 308 699 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=131490 $D=0
M1126 309 698 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=126860 $D=0
M1127 310 699 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=131490 $D=0
M1128 307 42 309 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=126860 $D=0
M1129 308 42 310 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=131490 $D=0
M1130 309 305 217 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=126860 $D=0
M1131 310 306 218 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=131490 $D=0
M1132 221 311 309 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=126860 $D=0
M1133 222 312 310 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=131490 $D=0
M1134 311 44 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=126860 $D=0
M1135 312 44 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=131490 $D=0
M1136 158 45 313 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=126860 $D=0
M1137 159 45 314 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=131490 $D=0
M1138 315 46 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=126860 $D=0
M1139 316 46 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=131490 $D=0
M1140 317 313 207 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=126860 $D=0
M1141 318 314 208 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=131490 $D=0
M1142 158 317 700 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=126860 $D=0
M1143 159 318 701 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=131490 $D=0
M1144 319 700 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=126860 $D=0
M1145 320 701 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=131490 $D=0
M1146 317 45 319 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=126860 $D=0
M1147 318 45 320 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=131490 $D=0
M1148 319 315 217 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=126860 $D=0
M1149 320 316 218 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=131490 $D=0
M1150 221 321 319 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=126860 $D=0
M1151 222 322 320 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=131490 $D=0
M1152 321 47 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=126860 $D=0
M1153 322 47 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=131490 $D=0
M1154 158 48 323 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=126860 $D=0
M1155 159 48 324 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=131490 $D=0
M1156 325 49 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=126860 $D=0
M1157 326 49 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=131490 $D=0
M1158 327 323 207 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=126860 $D=0
M1159 328 324 208 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=131490 $D=0
M1160 158 327 702 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=126860 $D=0
M1161 159 328 703 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=131490 $D=0
M1162 329 702 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=126860 $D=0
M1163 330 703 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=131490 $D=0
M1164 327 48 329 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=126860 $D=0
M1165 328 48 330 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=131490 $D=0
M1166 329 325 217 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=126860 $D=0
M1167 330 326 218 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=131490 $D=0
M1168 221 331 329 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=126860 $D=0
M1169 222 332 330 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=131490 $D=0
M1170 331 50 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=126860 $D=0
M1171 332 50 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=131490 $D=0
M1172 158 51 333 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=126860 $D=0
M1173 159 51 334 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=131490 $D=0
M1174 335 52 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=126860 $D=0
M1175 336 52 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=131490 $D=0
M1176 337 333 207 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=126860 $D=0
M1177 338 334 208 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=131490 $D=0
M1178 158 337 704 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=126860 $D=0
M1179 159 338 705 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=131490 $D=0
M1180 339 704 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=126860 $D=0
M1181 340 705 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=131490 $D=0
M1182 337 51 339 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=126860 $D=0
M1183 338 51 340 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=131490 $D=0
M1184 339 335 217 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=126860 $D=0
M1185 340 336 218 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=131490 $D=0
M1186 221 341 339 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=126860 $D=0
M1187 222 342 340 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=131490 $D=0
M1188 341 53 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=126860 $D=0
M1189 342 53 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=131490 $D=0
M1190 158 54 343 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=126860 $D=0
M1191 159 54 344 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=131490 $D=0
M1192 345 55 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=126860 $D=0
M1193 346 55 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=131490 $D=0
M1194 347 343 207 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=126860 $D=0
M1195 348 344 208 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=131490 $D=0
M1196 158 347 706 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=126860 $D=0
M1197 159 348 707 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=131490 $D=0
M1198 349 706 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=126860 $D=0
M1199 350 707 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=131490 $D=0
M1200 347 54 349 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=126860 $D=0
M1201 348 54 350 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=131490 $D=0
M1202 349 345 217 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=126860 $D=0
M1203 350 346 218 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=131490 $D=0
M1204 221 351 349 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=126860 $D=0
M1205 222 352 350 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=131490 $D=0
M1206 351 56 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=126860 $D=0
M1207 352 56 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=131490 $D=0
M1208 158 57 353 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=126860 $D=0
M1209 159 57 354 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=131490 $D=0
M1210 355 58 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=126860 $D=0
M1211 356 58 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=131490 $D=0
M1212 357 353 207 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=126860 $D=0
M1213 358 354 208 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=131490 $D=0
M1214 158 357 708 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=126860 $D=0
M1215 159 358 709 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=131490 $D=0
M1216 359 708 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=126860 $D=0
M1217 360 709 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=131490 $D=0
M1218 357 57 359 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=126860 $D=0
M1219 358 57 360 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=131490 $D=0
M1220 359 355 217 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=126860 $D=0
M1221 360 356 218 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=131490 $D=0
M1222 221 361 359 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=126860 $D=0
M1223 222 362 360 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=131490 $D=0
M1224 361 59 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=126860 $D=0
M1225 362 59 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=131490 $D=0
M1226 158 60 363 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=126860 $D=0
M1227 159 60 364 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=131490 $D=0
M1228 365 61 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=126860 $D=0
M1229 366 61 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=131490 $D=0
M1230 367 363 207 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=126860 $D=0
M1231 368 364 208 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=131490 $D=0
M1232 158 367 710 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=126860 $D=0
M1233 159 368 711 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=131490 $D=0
M1234 369 710 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=126860 $D=0
M1235 370 711 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=131490 $D=0
M1236 367 60 369 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=126860 $D=0
M1237 368 60 370 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=131490 $D=0
M1238 369 365 217 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=126860 $D=0
M1239 370 366 218 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=131490 $D=0
M1240 221 371 369 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=126860 $D=0
M1241 222 372 370 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=131490 $D=0
M1242 371 62 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=126860 $D=0
M1243 372 62 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=131490 $D=0
M1244 158 63 373 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=126860 $D=0
M1245 159 63 374 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=131490 $D=0
M1246 375 64 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=126860 $D=0
M1247 376 64 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=131490 $D=0
M1248 377 373 207 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=126860 $D=0
M1249 378 374 208 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=131490 $D=0
M1250 158 377 712 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=126860 $D=0
M1251 159 378 713 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=131490 $D=0
M1252 379 712 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=126860 $D=0
M1253 380 713 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=131490 $D=0
M1254 377 63 379 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=126860 $D=0
M1255 378 63 380 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=131490 $D=0
M1256 379 375 217 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=126860 $D=0
M1257 380 376 218 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=131490 $D=0
M1258 221 381 379 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=126860 $D=0
M1259 222 382 380 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=131490 $D=0
M1260 381 65 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=126860 $D=0
M1261 382 65 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=131490 $D=0
M1262 158 66 383 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=126860 $D=0
M1263 159 66 384 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=131490 $D=0
M1264 385 67 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=126860 $D=0
M1265 386 67 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=131490 $D=0
M1266 387 383 207 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=126860 $D=0
M1267 388 384 208 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=131490 $D=0
M1268 158 387 714 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=126860 $D=0
M1269 159 388 715 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=131490 $D=0
M1270 389 714 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=126860 $D=0
M1271 390 715 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=131490 $D=0
M1272 387 66 389 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=126860 $D=0
M1273 388 66 390 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=131490 $D=0
M1274 389 385 217 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=126860 $D=0
M1275 390 386 218 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=131490 $D=0
M1276 221 391 389 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=126860 $D=0
M1277 222 392 390 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=131490 $D=0
M1278 391 68 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=126860 $D=0
M1279 392 68 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=131490 $D=0
M1280 158 69 393 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=126860 $D=0
M1281 159 69 394 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=131490 $D=0
M1282 395 70 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=126860 $D=0
M1283 396 70 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=131490 $D=0
M1284 397 393 207 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=126860 $D=0
M1285 398 394 208 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=131490 $D=0
M1286 158 397 716 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=126860 $D=0
M1287 159 398 717 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=131490 $D=0
M1288 399 716 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=126860 $D=0
M1289 400 717 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=131490 $D=0
M1290 397 69 399 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=126860 $D=0
M1291 398 69 400 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=131490 $D=0
M1292 399 395 217 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=126860 $D=0
M1293 400 396 218 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=131490 $D=0
M1294 221 401 399 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=126860 $D=0
M1295 222 402 400 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=131490 $D=0
M1296 401 71 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=126860 $D=0
M1297 402 71 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=131490 $D=0
M1298 158 72 403 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=126860 $D=0
M1299 159 72 404 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=131490 $D=0
M1300 405 73 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=126860 $D=0
M1301 406 73 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=131490 $D=0
M1302 407 403 207 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=126860 $D=0
M1303 408 404 208 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=131490 $D=0
M1304 158 407 718 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=126860 $D=0
M1305 159 408 719 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=131490 $D=0
M1306 409 718 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=126860 $D=0
M1307 410 719 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=131490 $D=0
M1308 407 72 409 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=126860 $D=0
M1309 408 72 410 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=131490 $D=0
M1310 409 405 217 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=126860 $D=0
M1311 410 406 218 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=131490 $D=0
M1312 221 411 409 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=126860 $D=0
M1313 222 412 410 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=131490 $D=0
M1314 411 74 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=126860 $D=0
M1315 412 74 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=131490 $D=0
M1316 158 75 413 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=126860 $D=0
M1317 159 75 414 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=131490 $D=0
M1318 415 76 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=126860 $D=0
M1319 416 76 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=131490 $D=0
M1320 417 413 207 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=126860 $D=0
M1321 418 414 208 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=131490 $D=0
M1322 158 417 720 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=126860 $D=0
M1323 159 418 721 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=131490 $D=0
M1324 419 720 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=126860 $D=0
M1325 420 721 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=131490 $D=0
M1326 417 75 419 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=126860 $D=0
M1327 418 75 420 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=131490 $D=0
M1328 419 415 217 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=126860 $D=0
M1329 420 416 218 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=131490 $D=0
M1330 221 421 419 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=126860 $D=0
M1331 222 422 420 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=131490 $D=0
M1332 421 77 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=126860 $D=0
M1333 422 77 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=131490 $D=0
M1334 158 78 423 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=126860 $D=0
M1335 159 78 424 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=131490 $D=0
M1336 425 79 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=126860 $D=0
M1337 426 79 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=131490 $D=0
M1338 427 423 207 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=126860 $D=0
M1339 428 424 208 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=131490 $D=0
M1340 158 427 722 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=126860 $D=0
M1341 159 428 723 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=131490 $D=0
M1342 429 722 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=126860 $D=0
M1343 430 723 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=131490 $D=0
M1344 427 78 429 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=126860 $D=0
M1345 428 78 430 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=131490 $D=0
M1346 429 425 217 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=126860 $D=0
M1347 430 426 218 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=131490 $D=0
M1348 221 431 429 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=126860 $D=0
M1349 222 432 430 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=131490 $D=0
M1350 431 80 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=126860 $D=0
M1351 432 80 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=131490 $D=0
M1352 158 81 433 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=126860 $D=0
M1353 159 81 434 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=131490 $D=0
M1354 435 82 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=126860 $D=0
M1355 436 82 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=131490 $D=0
M1356 437 433 207 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=126860 $D=0
M1357 438 434 208 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=131490 $D=0
M1358 158 437 724 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=126860 $D=0
M1359 159 438 725 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=131490 $D=0
M1360 439 724 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=126860 $D=0
M1361 440 725 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=131490 $D=0
M1362 437 81 439 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=126860 $D=0
M1363 438 81 440 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=131490 $D=0
M1364 439 435 217 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=126860 $D=0
M1365 440 436 218 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=131490 $D=0
M1366 221 441 439 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=126860 $D=0
M1367 222 442 440 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=131490 $D=0
M1368 441 83 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=126860 $D=0
M1369 442 83 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=131490 $D=0
M1370 158 84 443 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=126860 $D=0
M1371 159 84 444 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=131490 $D=0
M1372 445 85 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=126860 $D=0
M1373 446 85 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=131490 $D=0
M1374 447 443 207 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=126860 $D=0
M1375 448 444 208 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=131490 $D=0
M1376 158 447 726 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=126860 $D=0
M1377 159 448 727 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=131490 $D=0
M1378 449 726 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=126860 $D=0
M1379 450 727 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=131490 $D=0
M1380 447 84 449 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=126860 $D=0
M1381 448 84 450 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=131490 $D=0
M1382 449 445 217 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=126860 $D=0
M1383 450 446 218 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=131490 $D=0
M1384 221 451 449 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=126860 $D=0
M1385 222 452 450 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=131490 $D=0
M1386 451 86 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=126860 $D=0
M1387 452 86 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=131490 $D=0
M1388 158 87 453 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=126860 $D=0
M1389 159 87 454 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=131490 $D=0
M1390 455 88 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=126860 $D=0
M1391 456 88 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=131490 $D=0
M1392 457 453 207 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=126860 $D=0
M1393 458 454 208 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=131490 $D=0
M1394 158 457 728 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=126860 $D=0
M1395 159 458 729 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=131490 $D=0
M1396 459 728 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=126860 $D=0
M1397 460 729 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=131490 $D=0
M1398 457 87 459 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=126860 $D=0
M1399 458 87 460 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=131490 $D=0
M1400 459 455 217 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=126860 $D=0
M1401 460 456 218 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=131490 $D=0
M1402 221 461 459 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=126860 $D=0
M1403 222 462 460 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=131490 $D=0
M1404 461 89 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=126860 $D=0
M1405 462 89 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=131490 $D=0
M1406 158 90 463 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=126860 $D=0
M1407 159 90 464 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=131490 $D=0
M1408 465 91 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=126860 $D=0
M1409 466 91 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=131490 $D=0
M1410 467 463 207 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=126860 $D=0
M1411 468 464 208 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=131490 $D=0
M1412 158 467 730 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=126860 $D=0
M1413 159 468 731 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=131490 $D=0
M1414 469 730 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=126860 $D=0
M1415 470 731 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=131490 $D=0
M1416 467 90 469 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=126860 $D=0
M1417 468 90 470 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=131490 $D=0
M1418 469 465 217 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=126860 $D=0
M1419 470 466 218 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=131490 $D=0
M1420 221 471 469 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=126860 $D=0
M1421 222 472 470 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=131490 $D=0
M1422 471 92 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=126860 $D=0
M1423 472 92 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=131490 $D=0
M1424 158 93 473 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=126860 $D=0
M1425 159 93 474 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=131490 $D=0
M1426 475 94 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=126860 $D=0
M1427 476 94 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=131490 $D=0
M1428 477 473 207 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=126860 $D=0
M1429 478 474 208 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=131490 $D=0
M1430 158 477 732 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=126860 $D=0
M1431 159 478 733 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=131490 $D=0
M1432 479 732 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=126860 $D=0
M1433 480 733 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=131490 $D=0
M1434 477 93 479 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=126860 $D=0
M1435 478 93 480 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=131490 $D=0
M1436 479 475 217 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=126860 $D=0
M1437 480 476 218 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=131490 $D=0
M1438 221 481 479 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=126860 $D=0
M1439 222 482 480 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=131490 $D=0
M1440 481 95 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=126860 $D=0
M1441 482 95 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=131490 $D=0
M1442 158 96 483 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=126860 $D=0
M1443 159 96 484 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=131490 $D=0
M1444 485 97 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=126860 $D=0
M1445 486 97 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=131490 $D=0
M1446 487 483 207 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=126860 $D=0
M1447 488 484 208 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=131490 $D=0
M1448 158 487 734 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=126860 $D=0
M1449 159 488 735 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=131490 $D=0
M1450 489 734 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=126860 $D=0
M1451 490 735 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=131490 $D=0
M1452 487 96 489 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=126860 $D=0
M1453 488 96 490 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=131490 $D=0
M1454 489 485 217 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=126860 $D=0
M1455 490 486 218 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=131490 $D=0
M1456 221 491 489 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=126860 $D=0
M1457 222 492 490 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=131490 $D=0
M1458 491 98 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=126860 $D=0
M1459 492 98 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=131490 $D=0
M1460 158 99 493 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=126860 $D=0
M1461 159 99 494 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=131490 $D=0
M1462 495 100 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=126860 $D=0
M1463 496 100 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=131490 $D=0
M1464 497 493 207 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=126860 $D=0
M1465 498 494 208 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=131490 $D=0
M1466 158 497 736 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=126860 $D=0
M1467 159 498 737 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=131490 $D=0
M1468 499 736 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=126860 $D=0
M1469 500 737 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=131490 $D=0
M1470 497 99 499 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=126860 $D=0
M1471 498 99 500 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=131490 $D=0
M1472 499 495 217 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=126860 $D=0
M1473 500 496 218 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=131490 $D=0
M1474 221 501 499 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=126860 $D=0
M1475 222 502 500 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=131490 $D=0
M1476 501 101 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=126860 $D=0
M1477 502 101 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=131490 $D=0
M1478 158 102 503 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=126860 $D=0
M1479 159 102 504 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=131490 $D=0
M1480 505 103 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=126860 $D=0
M1481 506 103 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=131490 $D=0
M1482 507 503 207 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=126860 $D=0
M1483 508 504 208 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=131490 $D=0
M1484 158 507 738 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=126860 $D=0
M1485 159 508 739 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=131490 $D=0
M1486 509 738 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=126860 $D=0
M1487 510 739 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=131490 $D=0
M1488 507 102 509 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=126860 $D=0
M1489 508 102 510 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=131490 $D=0
M1490 509 505 217 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=126860 $D=0
M1491 510 506 218 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=131490 $D=0
M1492 221 511 509 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=126860 $D=0
M1493 222 512 510 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=131490 $D=0
M1494 511 104 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=126860 $D=0
M1495 512 104 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=131490 $D=0
M1496 158 105 513 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=126860 $D=0
M1497 159 105 514 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=131490 $D=0
M1498 515 106 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=126860 $D=0
M1499 516 106 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=131490 $D=0
M1500 517 513 207 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=126860 $D=0
M1501 518 514 208 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=131490 $D=0
M1502 158 517 740 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=126860 $D=0
M1503 159 518 741 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=131490 $D=0
M1504 519 740 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=126860 $D=0
M1505 520 741 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=131490 $D=0
M1506 517 105 519 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=126860 $D=0
M1507 518 105 520 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=131490 $D=0
M1508 519 515 217 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=126860 $D=0
M1509 520 516 218 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=131490 $D=0
M1510 221 521 519 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=126860 $D=0
M1511 222 522 520 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=131490 $D=0
M1512 521 107 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=126860 $D=0
M1513 522 107 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=131490 $D=0
M1514 158 108 523 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=126860 $D=0
M1515 159 108 524 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=131490 $D=0
M1516 525 109 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=126860 $D=0
M1517 526 109 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=131490 $D=0
M1518 7 525 217 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=126860 $D=0
M1519 8 526 218 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=131490 $D=0
M1520 221 523 7 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=126860 $D=0
M1521 222 524 8 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=131490 $D=0
M1522 158 529 527 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=126860 $D=0
M1523 159 530 528 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=131490 $D=0
M1524 529 110 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=126860 $D=0
M1525 530 110 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=131490 $D=0
M1526 742 217 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=126860 $D=0
M1527 743 218 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=131490 $D=0
M1528 531 529 742 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=126860 $D=0
M1529 532 530 743 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=131490 $D=0
M1530 158 531 533 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=126860 $D=0
M1531 159 532 534 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=131490 $D=0
M1532 744 533 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=126860 $D=0
M1533 745 534 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=131490 $D=0
M1534 531 527 744 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=126860 $D=0
M1535 532 528 745 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=131490 $D=0
M1536 158 537 535 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=126860 $D=0
M1537 159 538 536 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=131490 $D=0
M1538 537 110 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=126860 $D=0
M1539 538 110 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=131490 $D=0
M1540 746 221 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=126860 $D=0
M1541 747 222 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=131490 $D=0
M1542 539 537 746 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=126860 $D=0
M1543 540 538 747 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=131490 $D=0
M1544 158 539 111 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=126860 $D=0
M1545 159 540 112 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=131490 $D=0
M1546 748 111 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=126860 $D=0
M1547 749 112 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=131490 $D=0
M1548 539 535 748 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=126860 $D=0
M1549 540 536 749 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=131490 $D=0
M1550 541 113 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=126860 $D=0
M1551 542 113 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=131490 $D=0
M1552 543 113 533 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=126860 $D=0
M1553 544 113 534 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=131490 $D=0
M1554 114 541 543 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=126860 $D=0
M1555 115 542 544 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=131490 $D=0
M1556 545 116 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=126860 $D=0
M1557 546 116 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=131490 $D=0
M1558 547 116 111 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=126860 $D=0
M1559 548 116 112 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=131490 $D=0
M1560 750 545 547 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=126860 $D=0
M1561 751 546 548 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=131490 $D=0
M1562 158 111 750 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=126860 $D=0
M1563 159 112 751 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=131490 $D=0
M1564 549 117 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=126860 $D=0
M1565 550 117 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=131490 $D=0
M1566 118 117 547 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=126860 $D=0
M1567 119 117 548 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=131490 $D=0
M1568 9 549 118 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=126860 $D=0
M1569 10 550 119 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=131490 $D=0
M1570 552 551 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=126860 $D=0
M1571 553 120 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=131490 $D=0
M1572 158 556 554 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=126860 $D=0
M1573 159 557 555 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=131490 $D=0
M1574 558 543 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=126860 $D=0
M1575 559 544 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=131490 $D=0
M1576 556 543 551 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=126860 $D=0
M1577 557 544 120 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=131490 $D=0
M1578 552 558 556 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=126860 $D=0
M1579 553 559 557 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=131490 $D=0
M1580 560 554 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=126860 $D=0
M1581 561 555 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=131490 $D=0
M1582 562 554 118 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=126860 $D=0
M1583 551 555 119 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=131490 $D=0
M1584 543 560 562 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=126860 $D=0
M1585 544 561 551 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=131490 $D=0
M1586 563 562 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=126860 $D=0
M1587 564 551 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=131490 $D=0
M1588 565 554 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=126860 $D=0
M1589 566 555 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=131490 $D=0
M1590 567 554 563 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=126860 $D=0
M1591 568 555 564 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=131490 $D=0
M1592 118 565 567 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=126860 $D=0
M1593 119 566 568 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=131490 $D=0
M1594 768 543 158 158 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=126500 $D=0
M1595 769 544 159 159 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=131130 $D=0
M1596 569 118 768 158 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=126500 $D=0
M1597 570 119 769 159 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=131130 $D=0
M1598 571 567 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=126860 $D=0
M1599 572 568 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=131490 $D=0
M1600 573 543 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=126860 $D=0
M1601 574 544 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=131490 $D=0
M1602 158 118 573 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=126860 $D=0
M1603 159 119 574 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=131490 $D=0
M1604 575 543 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=126860 $D=0
M1605 576 544 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=131490 $D=0
M1606 158 118 575 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=126860 $D=0
M1607 159 119 576 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=131490 $D=0
M1608 770 543 158 158 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=126680 $D=0
M1609 771 544 159 159 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=131310 $D=0
M1610 579 118 770 158 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=126680 $D=0
M1611 580 119 771 159 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=131310 $D=0
M1612 158 575 579 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=126860 $D=0
M1613 159 576 580 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=131490 $D=0
M1614 581 124 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=126860 $D=0
M1615 582 124 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=131490 $D=0
M1616 583 124 569 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=126860 $D=0
M1617 584 124 570 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=131490 $D=0
M1618 573 581 583 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=126860 $D=0
M1619 574 582 584 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=131490 $D=0
M1620 585 124 571 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=126860 $D=0
M1621 586 124 572 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=131490 $D=0
M1622 579 581 585 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=126860 $D=0
M1623 580 582 586 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=131490 $D=0
M1624 587 125 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=126860 $D=0
M1625 588 125 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=131490 $D=0
M1626 589 125 585 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=126860 $D=0
M1627 590 125 586 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=131490 $D=0
M1628 583 587 589 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=126860 $D=0
M1629 584 588 590 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=131490 $D=0
M1630 11 589 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=126860 $D=0
M1631 12 590 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=131490 $D=0
M1632 591 127 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=126860 $D=0
M1633 592 127 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=131490 $D=0
M1634 593 127 128 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=126860 $D=0
M1635 594 127 129 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=131490 $D=0
M1636 130 591 593 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=126860 $D=0
M1637 118 592 594 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=131490 $D=0
M1638 595 127 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=126860 $D=0
M1639 596 127 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=131490 $D=0
M1640 598 127 131 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=126860 $D=0
M1641 599 127 133 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=131490 $D=0
M1642 134 595 598 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=126860 $D=0
M1643 132 596 599 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=131490 $D=0
M1644 600 127 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=126860 $D=0
M1645 601 127 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=131490 $D=0
M1646 135 127 121 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=126860 $D=0
M1647 135 127 8 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=131490 $D=0
M1648 126 600 135 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=126860 $D=0
M1649 136 601 135 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=131490 $D=0
M1650 602 127 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=126860 $D=0
M1651 603 127 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=131490 $D=0
M1652 604 127 7 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=126860 $D=0
M1653 605 127 8 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=131490 $D=0
M1654 137 602 604 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=126860 $D=0
M1655 138 603 605 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=131490 $D=0
M1656 606 127 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=126860 $D=0
M1657 607 127 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=131490 $D=0
M1658 608 127 7 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=126860 $D=0
M1659 609 127 8 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=131490 $D=0
M1660 139 606 608 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=126860 $D=0
M1661 140 607 609 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=131490 $D=0
M1662 158 543 758 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=126860 $D=0
M1663 159 544 759 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=131490 $D=0
M1664 118 758 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=126860 $D=0
M1665 128 759 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=131490 $D=0
M1666 610 141 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=126860 $D=0
M1667 611 141 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=131490 $D=0
M1668 142 141 118 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=126860 $D=0
M1669 143 141 128 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=131490 $D=0
M1670 593 610 142 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=126860 $D=0
M1671 594 611 143 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=131490 $D=0
M1672 612 144 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=126860 $D=0
M1673 613 144 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=131490 $D=0
M1674 145 144 142 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=126860 $D=0
M1675 123 144 143 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=131490 $D=0
M1676 598 612 145 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=126860 $D=0
M1677 599 613 123 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=131490 $D=0
M1678 614 129 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=126860 $D=0
M1679 615 129 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=131490 $D=0
M1680 146 129 145 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=126860 $D=0
M1681 147 129 123 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=131490 $D=0
M1682 135 614 146 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=126860 $D=0
M1683 135 615 147 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=131490 $D=0
M1684 616 119 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=126860 $D=0
M1685 617 119 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=131490 $D=0
M1686 148 119 146 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=126860 $D=0
M1687 149 119 147 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=131490 $D=0
M1688 604 616 148 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=126860 $D=0
M1689 605 617 149 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=131490 $D=0
M1690 618 118 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=126860 $D=0
M1691 619 118 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=131490 $D=0
M1692 193 118 148 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=126860 $D=0
M1693 194 118 149 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=131490 $D=0
M1694 608 618 193 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=126860 $D=0
M1695 609 619 194 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=131490 $D=0
M1696 620 150 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=126860 $D=0
M1697 621 150 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=131490 $D=0
M1698 622 150 111 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=126860 $D=0
M1699 623 150 112 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=131490 $D=0
M1700 9 620 622 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=126860 $D=0
M1701 10 621 623 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=131490 $D=0
M1702 624 533 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=126860 $D=0
M1703 625 534 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=131490 $D=0
M1704 158 622 624 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=126860 $D=0
M1705 159 623 625 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=131490 $D=0
M1706 772 533 158 158 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=126680 $D=0
M1707 773 534 159 159 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=131310 $D=0
M1708 628 622 772 158 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=126680 $D=0
M1709 629 623 773 159 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=131310 $D=0
M1710 158 624 628 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=126860 $D=0
M1711 159 625 629 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=131490 $D=0
M1712 760 630 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=126860 $D=0
M1713 761 631 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=131490 $D=0
M1714 158 628 760 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=126860 $D=0
M1715 159 629 761 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=131490 $D=0
M1716 631 760 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=126860 $D=0
M1717 151 761 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=131490 $D=0
M1718 774 533 158 158 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=126500 $D=0
M1719 775 534 159 159 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=131130 $D=0
M1720 632 634 774 158 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=126500 $D=0
M1721 633 635 775 159 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=131130 $D=0
M1722 634 622 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=126860 $D=0
M1723 635 623 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=131490 $D=0
M1724 636 632 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=126860 $D=0
M1725 637 633 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=131490 $D=0
M1726 158 630 636 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=126860 $D=0
M1727 159 631 637 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=131490 $D=0
M1728 639 152 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=126860 $D=0
M1729 640 638 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=131490 $D=0
M1730 638 636 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=126860 $D=0
M1731 153 637 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=131490 $D=0
M1732 158 639 638 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=126860 $D=0
M1733 159 640 153 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=131490 $D=0
M1734 642 641 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=126860 $D=0
M1735 643 154 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=131490 $D=0
M1736 158 646 644 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=126860 $D=0
M1737 159 647 645 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=131490 $D=0
M1738 648 114 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=126860 $D=0
M1739 649 115 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=131490 $D=0
M1740 646 114 641 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=126860 $D=0
M1741 647 115 154 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=131490 $D=0
M1742 642 648 646 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=126860 $D=0
M1743 643 649 647 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=131490 $D=0
M1744 650 644 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=126860 $D=0
M1745 651 645 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=131490 $D=0
M1746 155 644 7 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=126860 $D=0
M1747 641 645 8 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=131490 $D=0
M1748 114 650 155 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=126860 $D=0
M1749 115 651 641 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=131490 $D=0
M1750 652 155 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=126860 $D=0
M1751 653 641 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=131490 $D=0
M1752 654 644 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=126860 $D=0
M1753 655 645 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=131490 $D=0
M1754 195 644 652 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=126860 $D=0
M1755 196 645 653 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=131490 $D=0
M1756 7 654 195 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=126860 $D=0
M1757 8 655 196 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=131490 $D=0
M1758 656 156 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=126860 $D=0
M1759 657 156 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=131490 $D=0
M1760 658 156 195 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=126860 $D=0
M1761 659 156 196 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=131490 $D=0
M1762 11 656 658 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=126860 $D=0
M1763 12 657 659 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=131490 $D=0
M1764 660 157 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=126860 $D=0
M1765 661 157 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=131490 $D=0
M1766 157 157 658 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=126860 $D=0
M1767 157 157 659 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=131490 $D=0
M1768 7 660 157 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=126860 $D=0
M1769 8 661 157 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=131490 $D=0
M1770 662 110 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=126860 $D=0
M1771 663 110 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=131490 $D=0
M1772 158 662 664 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=126860 $D=0
M1773 159 663 665 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=131490 $D=0
M1774 666 110 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=126860 $D=0
M1775 667 110 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=131490 $D=0
M1776 668 664 157 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=126860 $D=0
M1777 669 665 157 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=131490 $D=0
M1778 158 668 762 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=126860 $D=0
M1779 159 669 763 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=131490 $D=0
M1780 670 762 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=126860 $D=0
M1781 671 763 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=131490 $D=0
M1782 668 662 670 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=126860 $D=0
M1783 669 663 671 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=131490 $D=0
M1784 672 666 670 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=126860 $D=0
M1785 673 667 671 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=131490 $D=0
M1786 158 676 674 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=126860 $D=0
M1787 159 677 675 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=131490 $D=0
M1788 676 110 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=126860 $D=0
M1789 677 110 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=131490 $D=0
M1790 764 672 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=126860 $D=0
M1791 765 673 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=131490 $D=0
M1792 678 676 764 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=126860 $D=0
M1793 679 677 765 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=131490 $D=0
M1794 158 678 114 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=126860 $D=0
M1795 159 679 115 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=131490 $D=0
M1796 766 114 158 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=126860 $D=0
M1797 767 115 159 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=131490 $D=0
M1798 678 674 766 158 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=126860 $D=0
M1799 679 675 767 159 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=131490 $D=0
.ENDS
***************************************
.SUBCKT ICV_26 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141
+ 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161
+ 162
** N=800 EP=161 IP=1514 FDC=1800
M0 175 1 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=116350 $D=1
M1 176 1 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=120980 $D=1
M2 177 175 2 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=116350 $D=1
M3 178 176 3 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=120980 $D=1
M4 7 1 177 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=116350 $D=1
M5 8 1 178 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=120980 $D=1
M6 179 175 2 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=116350 $D=1
M7 180 176 3 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=120980 $D=1
M8 2 1 179 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=116350 $D=1
M9 3 1 180 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=120980 $D=1
M10 181 175 2 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=116350 $D=1
M11 182 176 3 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=120980 $D=1
M12 2 1 181 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=116350 $D=1
M13 3 1 182 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=120980 $D=1
M14 185 183 181 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=116350 $D=1
M15 186 184 182 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=120980 $D=1
M16 183 4 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=116350 $D=1
M17 184 4 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=120980 $D=1
M18 187 183 179 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=116350 $D=1
M19 188 184 180 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=120980 $D=1
M20 177 4 187 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=116350 $D=1
M21 178 4 188 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=120980 $D=1
M22 189 5 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=116350 $D=1
M23 190 5 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=120980 $D=1
M24 191 189 187 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=116350 $D=1
M25 192 190 188 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=120980 $D=1
M26 185 5 191 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=116350 $D=1
M27 186 5 192 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=120980 $D=1
M28 193 6 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=116350 $D=1
M29 194 6 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=120980 $D=1
M30 195 193 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=116350 $D=1
M31 196 194 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=120980 $D=1
M32 9 6 195 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=116350 $D=1
M33 10 6 196 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=120980 $D=1
M34 197 193 11 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=116350 $D=1
M35 198 194 12 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=120980 $D=1
M36 199 6 197 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=116350 $D=1
M37 200 6 198 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=120980 $D=1
M38 203 193 201 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=116350 $D=1
M39 204 194 202 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=120980 $D=1
M40 191 6 203 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=116350 $D=1
M41 192 6 204 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=120980 $D=1
M42 207 205 203 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=116350 $D=1
M43 208 206 204 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=120980 $D=1
M44 205 13 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=116350 $D=1
M45 206 13 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=120980 $D=1
M46 209 205 197 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=116350 $D=1
M47 210 206 198 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=120980 $D=1
M48 195 13 209 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=116350 $D=1
M49 196 13 210 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=120980 $D=1
M50 211 14 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=116350 $D=1
M51 212 14 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=120980 $D=1
M52 213 211 209 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=116350 $D=1
M53 214 212 210 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=120980 $D=1
M54 207 14 213 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=116350 $D=1
M55 208 14 214 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=120980 $D=1
M56 7 15 215 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=116350 $D=1
M57 8 15 216 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=120980 $D=1
M58 217 16 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=116350 $D=1
M59 218 16 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=120980 $D=1
M60 219 15 213 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=116350 $D=1
M61 220 15 214 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=120980 $D=1
M62 7 219 689 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=116350 $D=1
M63 8 220 690 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=120980 $D=1
M64 221 689 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=116350 $D=1
M65 222 690 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=120980 $D=1
M66 219 215 221 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=116350 $D=1
M67 220 216 222 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=120980 $D=1
M68 221 16 223 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=116350 $D=1
M69 222 16 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=120980 $D=1
M70 227 17 221 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=116350 $D=1
M71 228 17 222 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=120980 $D=1
M72 225 17 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=116350 $D=1
M73 226 17 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=120980 $D=1
M74 7 18 229 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=116350 $D=1
M75 8 18 230 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=120980 $D=1
M76 231 19 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=116350 $D=1
M77 232 19 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=120980 $D=1
M78 233 18 213 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=116350 $D=1
M79 234 18 214 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=120980 $D=1
M80 7 233 691 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=116350 $D=1
M81 8 234 692 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=120980 $D=1
M82 235 691 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=116350 $D=1
M83 236 692 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=120980 $D=1
M84 233 229 235 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=116350 $D=1
M85 234 230 236 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=120980 $D=1
M86 235 19 223 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=116350 $D=1
M87 236 19 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=120980 $D=1
M88 227 20 235 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=116350 $D=1
M89 228 20 236 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=120980 $D=1
M90 237 20 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=116350 $D=1
M91 238 20 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=120980 $D=1
M92 7 21 239 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=116350 $D=1
M93 8 21 240 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=120980 $D=1
M94 241 22 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=116350 $D=1
M95 242 22 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=120980 $D=1
M96 243 21 213 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=116350 $D=1
M97 244 21 214 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=120980 $D=1
M98 7 243 693 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=116350 $D=1
M99 8 244 694 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=120980 $D=1
M100 245 693 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=116350 $D=1
M101 246 694 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=120980 $D=1
M102 243 239 245 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=116350 $D=1
M103 244 240 246 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=120980 $D=1
M104 245 22 223 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=116350 $D=1
M105 246 22 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=120980 $D=1
M106 227 23 245 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=116350 $D=1
M107 228 23 246 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=120980 $D=1
M108 247 23 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=116350 $D=1
M109 248 23 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=120980 $D=1
M110 7 24 249 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=116350 $D=1
M111 8 24 250 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=120980 $D=1
M112 251 25 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=116350 $D=1
M113 252 25 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=120980 $D=1
M114 253 24 213 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=116350 $D=1
M115 254 24 214 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=120980 $D=1
M116 7 253 695 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=116350 $D=1
M117 8 254 696 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=120980 $D=1
M118 255 695 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=116350 $D=1
M119 256 696 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=120980 $D=1
M120 253 249 255 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=116350 $D=1
M121 254 250 256 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=120980 $D=1
M122 255 25 223 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=116350 $D=1
M123 256 25 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=120980 $D=1
M124 227 26 255 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=116350 $D=1
M125 228 26 256 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=120980 $D=1
M126 257 26 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=116350 $D=1
M127 258 26 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=120980 $D=1
M128 7 27 259 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=116350 $D=1
M129 8 27 260 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=120980 $D=1
M130 261 28 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=116350 $D=1
M131 262 28 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=120980 $D=1
M132 263 27 213 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=116350 $D=1
M133 264 27 214 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=120980 $D=1
M134 7 263 697 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=116350 $D=1
M135 8 264 698 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=120980 $D=1
M136 265 697 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=116350 $D=1
M137 266 698 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=120980 $D=1
M138 263 259 265 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=116350 $D=1
M139 264 260 266 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=120980 $D=1
M140 265 28 223 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=116350 $D=1
M141 266 28 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=120980 $D=1
M142 227 29 265 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=116350 $D=1
M143 228 29 266 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=120980 $D=1
M144 267 29 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=116350 $D=1
M145 268 29 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=120980 $D=1
M146 7 30 269 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=116350 $D=1
M147 8 30 270 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=120980 $D=1
M148 271 31 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=116350 $D=1
M149 272 31 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=120980 $D=1
M150 273 30 213 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=116350 $D=1
M151 274 30 214 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=120980 $D=1
M152 7 273 699 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=116350 $D=1
M153 8 274 700 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=120980 $D=1
M154 275 699 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=116350 $D=1
M155 276 700 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=120980 $D=1
M156 273 269 275 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=116350 $D=1
M157 274 270 276 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=120980 $D=1
M158 275 31 223 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=116350 $D=1
M159 276 31 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=120980 $D=1
M160 227 32 275 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=116350 $D=1
M161 228 32 276 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=120980 $D=1
M162 277 32 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=116350 $D=1
M163 278 32 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=120980 $D=1
M164 7 33 279 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=116350 $D=1
M165 8 33 280 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=120980 $D=1
M166 281 34 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=116350 $D=1
M167 282 34 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=120980 $D=1
M168 283 33 213 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=116350 $D=1
M169 284 33 214 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=120980 $D=1
M170 7 283 701 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=116350 $D=1
M171 8 284 702 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=120980 $D=1
M172 285 701 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=116350 $D=1
M173 286 702 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=120980 $D=1
M174 283 279 285 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=116350 $D=1
M175 284 280 286 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=120980 $D=1
M176 285 34 223 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=116350 $D=1
M177 286 34 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=120980 $D=1
M178 227 35 285 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=116350 $D=1
M179 228 35 286 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=120980 $D=1
M180 287 35 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=116350 $D=1
M181 288 35 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=120980 $D=1
M182 7 36 289 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=116350 $D=1
M183 8 36 290 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=120980 $D=1
M184 291 37 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=116350 $D=1
M185 292 37 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=120980 $D=1
M186 293 36 213 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=116350 $D=1
M187 294 36 214 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=120980 $D=1
M188 7 293 703 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=116350 $D=1
M189 8 294 704 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=120980 $D=1
M190 295 703 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=116350 $D=1
M191 296 704 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=120980 $D=1
M192 293 289 295 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=116350 $D=1
M193 294 290 296 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=120980 $D=1
M194 295 37 223 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=116350 $D=1
M195 296 37 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=120980 $D=1
M196 227 38 295 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=116350 $D=1
M197 228 38 296 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=120980 $D=1
M198 297 38 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=116350 $D=1
M199 298 38 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=120980 $D=1
M200 7 39 299 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=116350 $D=1
M201 8 39 300 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=120980 $D=1
M202 301 40 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=116350 $D=1
M203 302 40 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=120980 $D=1
M204 303 39 213 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=116350 $D=1
M205 304 39 214 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=120980 $D=1
M206 7 303 705 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=116350 $D=1
M207 8 304 706 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=120980 $D=1
M208 305 705 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=116350 $D=1
M209 306 706 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=120980 $D=1
M210 303 299 305 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=116350 $D=1
M211 304 300 306 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=120980 $D=1
M212 305 40 223 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=116350 $D=1
M213 306 40 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=120980 $D=1
M214 227 41 305 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=116350 $D=1
M215 228 41 306 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=120980 $D=1
M216 307 41 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=116350 $D=1
M217 308 41 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=120980 $D=1
M218 7 42 309 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=116350 $D=1
M219 8 42 310 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=120980 $D=1
M220 311 43 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=116350 $D=1
M221 312 43 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=120980 $D=1
M222 313 42 213 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=116350 $D=1
M223 314 42 214 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=120980 $D=1
M224 7 313 707 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=116350 $D=1
M225 8 314 708 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=120980 $D=1
M226 315 707 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=116350 $D=1
M227 316 708 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=120980 $D=1
M228 313 309 315 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=116350 $D=1
M229 314 310 316 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=120980 $D=1
M230 315 43 223 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=116350 $D=1
M231 316 43 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=120980 $D=1
M232 227 44 315 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=116350 $D=1
M233 228 44 316 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=120980 $D=1
M234 317 44 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=116350 $D=1
M235 318 44 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=120980 $D=1
M236 7 45 319 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=116350 $D=1
M237 8 45 320 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=120980 $D=1
M238 321 46 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=116350 $D=1
M239 322 46 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=120980 $D=1
M240 323 45 213 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=116350 $D=1
M241 324 45 214 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=120980 $D=1
M242 7 323 709 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=116350 $D=1
M243 8 324 710 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=120980 $D=1
M244 325 709 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=116350 $D=1
M245 326 710 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=120980 $D=1
M246 323 319 325 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=116350 $D=1
M247 324 320 326 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=120980 $D=1
M248 325 46 223 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=116350 $D=1
M249 326 46 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=120980 $D=1
M250 227 47 325 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=116350 $D=1
M251 228 47 326 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=120980 $D=1
M252 327 47 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=116350 $D=1
M253 328 47 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=120980 $D=1
M254 7 48 329 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=116350 $D=1
M255 8 48 330 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=120980 $D=1
M256 331 49 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=116350 $D=1
M257 332 49 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=120980 $D=1
M258 333 48 213 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=116350 $D=1
M259 334 48 214 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=120980 $D=1
M260 7 333 711 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=116350 $D=1
M261 8 334 712 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=120980 $D=1
M262 335 711 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=116350 $D=1
M263 336 712 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=120980 $D=1
M264 333 329 335 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=116350 $D=1
M265 334 330 336 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=120980 $D=1
M266 335 49 223 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=116350 $D=1
M267 336 49 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=120980 $D=1
M268 227 50 335 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=116350 $D=1
M269 228 50 336 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=120980 $D=1
M270 337 50 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=116350 $D=1
M271 338 50 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=120980 $D=1
M272 7 51 339 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=116350 $D=1
M273 8 51 340 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=120980 $D=1
M274 341 52 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=116350 $D=1
M275 342 52 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=120980 $D=1
M276 343 51 213 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=116350 $D=1
M277 344 51 214 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=120980 $D=1
M278 7 343 713 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=116350 $D=1
M279 8 344 714 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=120980 $D=1
M280 345 713 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=116350 $D=1
M281 346 714 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=120980 $D=1
M282 343 339 345 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=116350 $D=1
M283 344 340 346 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=120980 $D=1
M284 345 52 223 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=116350 $D=1
M285 346 52 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=120980 $D=1
M286 227 53 345 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=116350 $D=1
M287 228 53 346 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=120980 $D=1
M288 347 53 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=116350 $D=1
M289 348 53 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=120980 $D=1
M290 7 54 349 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=116350 $D=1
M291 8 54 350 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=120980 $D=1
M292 351 55 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=116350 $D=1
M293 352 55 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=120980 $D=1
M294 353 54 213 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=116350 $D=1
M295 354 54 214 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=120980 $D=1
M296 7 353 715 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=116350 $D=1
M297 8 354 716 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=120980 $D=1
M298 355 715 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=116350 $D=1
M299 356 716 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=120980 $D=1
M300 353 349 355 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=116350 $D=1
M301 354 350 356 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=120980 $D=1
M302 355 55 223 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=116350 $D=1
M303 356 55 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=120980 $D=1
M304 227 56 355 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=116350 $D=1
M305 228 56 356 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=120980 $D=1
M306 357 56 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=116350 $D=1
M307 358 56 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=120980 $D=1
M308 7 57 359 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=116350 $D=1
M309 8 57 360 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=120980 $D=1
M310 361 58 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=116350 $D=1
M311 362 58 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=120980 $D=1
M312 363 57 213 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=116350 $D=1
M313 364 57 214 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=120980 $D=1
M314 7 363 717 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=116350 $D=1
M315 8 364 718 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=120980 $D=1
M316 365 717 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=116350 $D=1
M317 366 718 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=120980 $D=1
M318 363 359 365 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=116350 $D=1
M319 364 360 366 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=120980 $D=1
M320 365 58 223 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=116350 $D=1
M321 366 58 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=120980 $D=1
M322 227 59 365 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=116350 $D=1
M323 228 59 366 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=120980 $D=1
M324 367 59 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=116350 $D=1
M325 368 59 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=120980 $D=1
M326 7 60 369 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=116350 $D=1
M327 8 60 370 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=120980 $D=1
M328 371 61 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=116350 $D=1
M329 372 61 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=120980 $D=1
M330 373 60 213 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=116350 $D=1
M331 374 60 214 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=120980 $D=1
M332 7 373 719 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=116350 $D=1
M333 8 374 720 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=120980 $D=1
M334 375 719 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=116350 $D=1
M335 376 720 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=120980 $D=1
M336 373 369 375 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=116350 $D=1
M337 374 370 376 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=120980 $D=1
M338 375 61 223 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=116350 $D=1
M339 376 61 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=120980 $D=1
M340 227 62 375 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=116350 $D=1
M341 228 62 376 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=120980 $D=1
M342 377 62 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=116350 $D=1
M343 378 62 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=120980 $D=1
M344 7 63 379 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=116350 $D=1
M345 8 63 380 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=120980 $D=1
M346 381 64 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=116350 $D=1
M347 382 64 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=120980 $D=1
M348 383 63 213 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=116350 $D=1
M349 384 63 214 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=120980 $D=1
M350 7 383 721 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=116350 $D=1
M351 8 384 722 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=120980 $D=1
M352 385 721 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=116350 $D=1
M353 386 722 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=120980 $D=1
M354 383 379 385 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=116350 $D=1
M355 384 380 386 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=120980 $D=1
M356 385 64 223 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=116350 $D=1
M357 386 64 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=120980 $D=1
M358 227 65 385 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=116350 $D=1
M359 228 65 386 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=120980 $D=1
M360 387 65 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=116350 $D=1
M361 388 65 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=120980 $D=1
M362 7 66 389 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=116350 $D=1
M363 8 66 390 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=120980 $D=1
M364 391 67 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=116350 $D=1
M365 392 67 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=120980 $D=1
M366 393 66 213 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=116350 $D=1
M367 394 66 214 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=120980 $D=1
M368 7 393 723 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=116350 $D=1
M369 8 394 724 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=120980 $D=1
M370 395 723 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=116350 $D=1
M371 396 724 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=120980 $D=1
M372 393 389 395 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=116350 $D=1
M373 394 390 396 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=120980 $D=1
M374 395 67 223 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=116350 $D=1
M375 396 67 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=120980 $D=1
M376 227 68 395 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=116350 $D=1
M377 228 68 396 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=120980 $D=1
M378 397 68 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=116350 $D=1
M379 398 68 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=120980 $D=1
M380 7 69 399 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=116350 $D=1
M381 8 69 400 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=120980 $D=1
M382 401 70 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=116350 $D=1
M383 402 70 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=120980 $D=1
M384 403 69 213 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=116350 $D=1
M385 404 69 214 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=120980 $D=1
M386 7 403 725 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=116350 $D=1
M387 8 404 726 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=120980 $D=1
M388 405 725 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=116350 $D=1
M389 406 726 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=120980 $D=1
M390 403 399 405 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=116350 $D=1
M391 404 400 406 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=120980 $D=1
M392 405 70 223 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=116350 $D=1
M393 406 70 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=120980 $D=1
M394 227 71 405 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=116350 $D=1
M395 228 71 406 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=120980 $D=1
M396 407 71 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=116350 $D=1
M397 408 71 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=120980 $D=1
M398 7 72 409 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=116350 $D=1
M399 8 72 410 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=120980 $D=1
M400 411 73 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=116350 $D=1
M401 412 73 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=120980 $D=1
M402 413 72 213 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=116350 $D=1
M403 414 72 214 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=120980 $D=1
M404 7 413 727 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=116350 $D=1
M405 8 414 728 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=120980 $D=1
M406 415 727 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=116350 $D=1
M407 416 728 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=120980 $D=1
M408 413 409 415 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=116350 $D=1
M409 414 410 416 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=120980 $D=1
M410 415 73 223 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=116350 $D=1
M411 416 73 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=120980 $D=1
M412 227 74 415 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=116350 $D=1
M413 228 74 416 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=120980 $D=1
M414 417 74 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=116350 $D=1
M415 418 74 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=120980 $D=1
M416 7 75 419 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=116350 $D=1
M417 8 75 420 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=120980 $D=1
M418 421 76 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=116350 $D=1
M419 422 76 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=120980 $D=1
M420 423 75 213 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=116350 $D=1
M421 424 75 214 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=120980 $D=1
M422 7 423 729 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=116350 $D=1
M423 8 424 730 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=120980 $D=1
M424 425 729 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=116350 $D=1
M425 426 730 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=120980 $D=1
M426 423 419 425 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=116350 $D=1
M427 424 420 426 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=120980 $D=1
M428 425 76 223 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=116350 $D=1
M429 426 76 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=120980 $D=1
M430 227 77 425 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=116350 $D=1
M431 228 77 426 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=120980 $D=1
M432 427 77 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=116350 $D=1
M433 428 77 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=120980 $D=1
M434 7 78 429 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=116350 $D=1
M435 8 78 430 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=120980 $D=1
M436 431 79 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=116350 $D=1
M437 432 79 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=120980 $D=1
M438 433 78 213 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=116350 $D=1
M439 434 78 214 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=120980 $D=1
M440 7 433 731 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=116350 $D=1
M441 8 434 732 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=120980 $D=1
M442 435 731 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=116350 $D=1
M443 436 732 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=120980 $D=1
M444 433 429 435 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=116350 $D=1
M445 434 430 436 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=120980 $D=1
M446 435 79 223 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=116350 $D=1
M447 436 79 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=120980 $D=1
M448 227 80 435 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=116350 $D=1
M449 228 80 436 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=120980 $D=1
M450 437 80 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=116350 $D=1
M451 438 80 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=120980 $D=1
M452 7 81 439 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=116350 $D=1
M453 8 81 440 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=120980 $D=1
M454 441 82 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=116350 $D=1
M455 442 82 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=120980 $D=1
M456 443 81 213 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=116350 $D=1
M457 444 81 214 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=120980 $D=1
M458 7 443 733 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=116350 $D=1
M459 8 444 734 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=120980 $D=1
M460 445 733 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=116350 $D=1
M461 446 734 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=120980 $D=1
M462 443 439 445 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=116350 $D=1
M463 444 440 446 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=120980 $D=1
M464 445 82 223 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=116350 $D=1
M465 446 82 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=120980 $D=1
M466 227 83 445 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=116350 $D=1
M467 228 83 446 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=120980 $D=1
M468 447 83 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=116350 $D=1
M469 448 83 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=120980 $D=1
M470 7 84 449 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=116350 $D=1
M471 8 84 450 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=120980 $D=1
M472 451 85 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=116350 $D=1
M473 452 85 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=120980 $D=1
M474 453 84 213 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=116350 $D=1
M475 454 84 214 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=120980 $D=1
M476 7 453 735 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=116350 $D=1
M477 8 454 736 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=120980 $D=1
M478 455 735 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=116350 $D=1
M479 456 736 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=120980 $D=1
M480 453 449 455 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=116350 $D=1
M481 454 450 456 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=120980 $D=1
M482 455 85 223 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=116350 $D=1
M483 456 85 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=120980 $D=1
M484 227 86 455 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=116350 $D=1
M485 228 86 456 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=120980 $D=1
M486 457 86 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=116350 $D=1
M487 458 86 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=120980 $D=1
M488 7 87 459 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=116350 $D=1
M489 8 87 460 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=120980 $D=1
M490 461 88 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=116350 $D=1
M491 462 88 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=120980 $D=1
M492 463 87 213 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=116350 $D=1
M493 464 87 214 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=120980 $D=1
M494 7 463 737 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=116350 $D=1
M495 8 464 738 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=120980 $D=1
M496 465 737 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=116350 $D=1
M497 466 738 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=120980 $D=1
M498 463 459 465 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=116350 $D=1
M499 464 460 466 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=120980 $D=1
M500 465 88 223 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=116350 $D=1
M501 466 88 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=120980 $D=1
M502 227 89 465 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=116350 $D=1
M503 228 89 466 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=120980 $D=1
M504 467 89 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=116350 $D=1
M505 468 89 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=120980 $D=1
M506 7 90 469 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=116350 $D=1
M507 8 90 470 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=120980 $D=1
M508 471 91 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=116350 $D=1
M509 472 91 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=120980 $D=1
M510 473 90 213 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=116350 $D=1
M511 474 90 214 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=120980 $D=1
M512 7 473 739 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=116350 $D=1
M513 8 474 740 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=120980 $D=1
M514 475 739 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=116350 $D=1
M515 476 740 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=120980 $D=1
M516 473 469 475 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=116350 $D=1
M517 474 470 476 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=120980 $D=1
M518 475 91 223 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=116350 $D=1
M519 476 91 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=120980 $D=1
M520 227 92 475 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=116350 $D=1
M521 228 92 476 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=120980 $D=1
M522 477 92 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=116350 $D=1
M523 478 92 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=120980 $D=1
M524 7 93 479 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=116350 $D=1
M525 8 93 480 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=120980 $D=1
M526 481 94 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=116350 $D=1
M527 482 94 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=120980 $D=1
M528 483 93 213 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=116350 $D=1
M529 484 93 214 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=120980 $D=1
M530 7 483 741 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=116350 $D=1
M531 8 484 742 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=120980 $D=1
M532 485 741 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=116350 $D=1
M533 486 742 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=120980 $D=1
M534 483 479 485 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=116350 $D=1
M535 484 480 486 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=120980 $D=1
M536 485 94 223 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=116350 $D=1
M537 486 94 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=120980 $D=1
M538 227 95 485 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=116350 $D=1
M539 228 95 486 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=120980 $D=1
M540 487 95 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=116350 $D=1
M541 488 95 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=120980 $D=1
M542 7 96 489 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=116350 $D=1
M543 8 96 490 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=120980 $D=1
M544 491 97 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=116350 $D=1
M545 492 97 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=120980 $D=1
M546 493 96 213 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=116350 $D=1
M547 494 96 214 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=120980 $D=1
M548 7 493 743 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=116350 $D=1
M549 8 494 744 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=120980 $D=1
M550 495 743 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=116350 $D=1
M551 496 744 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=120980 $D=1
M552 493 489 495 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=116350 $D=1
M553 494 490 496 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=120980 $D=1
M554 495 97 223 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=116350 $D=1
M555 496 97 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=120980 $D=1
M556 227 98 495 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=116350 $D=1
M557 228 98 496 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=120980 $D=1
M558 497 98 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=116350 $D=1
M559 498 98 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=120980 $D=1
M560 7 99 499 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=116350 $D=1
M561 8 99 500 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=120980 $D=1
M562 501 100 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=116350 $D=1
M563 502 100 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=120980 $D=1
M564 503 99 213 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=116350 $D=1
M565 504 99 214 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=120980 $D=1
M566 7 503 745 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=116350 $D=1
M567 8 504 746 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=120980 $D=1
M568 505 745 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=116350 $D=1
M569 506 746 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=120980 $D=1
M570 503 499 505 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=116350 $D=1
M571 504 500 506 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=120980 $D=1
M572 505 100 223 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=116350 $D=1
M573 506 100 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=120980 $D=1
M574 227 101 505 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=116350 $D=1
M575 228 101 506 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=120980 $D=1
M576 507 101 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=116350 $D=1
M577 508 101 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=120980 $D=1
M578 7 102 509 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=116350 $D=1
M579 8 102 510 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=120980 $D=1
M580 511 103 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=116350 $D=1
M581 512 103 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=120980 $D=1
M582 513 102 213 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=116350 $D=1
M583 514 102 214 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=120980 $D=1
M584 7 513 747 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=116350 $D=1
M585 8 514 748 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=120980 $D=1
M586 515 747 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=116350 $D=1
M587 516 748 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=120980 $D=1
M588 513 509 515 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=116350 $D=1
M589 514 510 516 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=120980 $D=1
M590 515 103 223 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=116350 $D=1
M591 516 103 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=120980 $D=1
M592 227 104 515 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=116350 $D=1
M593 228 104 516 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=120980 $D=1
M594 517 104 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=116350 $D=1
M595 518 104 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=120980 $D=1
M596 7 105 519 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=116350 $D=1
M597 8 105 520 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=120980 $D=1
M598 521 106 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=116350 $D=1
M599 522 106 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=120980 $D=1
M600 523 105 213 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=116350 $D=1
M601 524 105 214 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=120980 $D=1
M602 7 523 749 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=116350 $D=1
M603 8 524 750 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=120980 $D=1
M604 525 749 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=116350 $D=1
M605 526 750 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=120980 $D=1
M606 523 519 525 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=116350 $D=1
M607 524 520 526 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=120980 $D=1
M608 525 106 223 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=116350 $D=1
M609 526 106 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=120980 $D=1
M610 227 107 525 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=116350 $D=1
M611 228 107 526 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=120980 $D=1
M612 527 107 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=116350 $D=1
M613 528 107 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=120980 $D=1
M614 7 108 529 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=116350 $D=1
M615 8 108 530 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=120980 $D=1
M616 531 109 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=116350 $D=1
M617 532 109 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=120980 $D=1
M618 7 109 223 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=116350 $D=1
M619 8 109 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=120980 $D=1
M620 227 108 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=116350 $D=1
M621 228 108 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=120980 $D=1
M622 7 535 533 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=116350 $D=1
M623 8 536 534 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=120980 $D=1
M624 535 110 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=116350 $D=1
M625 536 110 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=120980 $D=1
M626 751 223 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=116350 $D=1
M627 752 224 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=120980 $D=1
M628 537 533 751 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=116350 $D=1
M629 538 534 752 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=120980 $D=1
M630 7 537 539 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=116350 $D=1
M631 8 538 540 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=120980 $D=1
M632 753 539 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=116350 $D=1
M633 754 540 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=120980 $D=1
M634 537 535 753 7 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=116350 $D=1
M635 538 536 754 8 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=120980 $D=1
M636 7 543 541 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=116350 $D=1
M637 8 544 542 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=120980 $D=1
M638 543 110 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=116350 $D=1
M639 544 110 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=120980 $D=1
M640 755 227 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=116350 $D=1
M641 756 228 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=120980 $D=1
M642 545 541 755 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=116350 $D=1
M643 546 542 756 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=120980 $D=1
M644 7 545 111 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=116350 $D=1
M645 8 546 112 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=120980 $D=1
M646 757 111 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=116350 $D=1
M647 758 112 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=120980 $D=1
M648 545 543 757 7 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=116350 $D=1
M649 546 544 758 8 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=120980 $D=1
M650 547 113 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=116350 $D=1
M651 548 113 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=120980 $D=1
M652 549 547 539 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=116350 $D=1
M653 550 548 540 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=120980 $D=1
M654 114 113 549 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=116350 $D=1
M655 115 113 550 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=120980 $D=1
M656 551 116 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=116350 $D=1
M657 552 116 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=120980 $D=1
M658 553 551 111 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=116350 $D=1
M659 554 552 112 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=120980 $D=1
M660 759 116 553 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=116350 $D=1
M661 760 116 554 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=120980 $D=1
M662 7 111 759 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=116350 $D=1
M663 8 112 760 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=120980 $D=1
M664 555 117 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=116350 $D=1
M665 556 117 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=120980 $D=1
M666 557 555 553 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=116350 $D=1
M667 558 556 554 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=120980 $D=1
M668 9 117 557 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=116350 $D=1
M669 10 117 558 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=120980 $D=1
M670 560 559 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=116350 $D=1
M671 561 118 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=120980 $D=1
M672 7 564 562 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=116350 $D=1
M673 8 565 563 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=120980 $D=1
M674 566 549 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=116350 $D=1
M675 567 550 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=120980 $D=1
M676 564 566 559 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=116350 $D=1
M677 565 567 118 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=120980 $D=1
M678 560 549 564 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=116350 $D=1
M679 561 550 565 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=120980 $D=1
M680 568 562 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=116350 $D=1
M681 569 563 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=120980 $D=1
M682 119 568 557 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=116350 $D=1
M683 559 569 558 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=120980 $D=1
M684 549 562 119 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=116350 $D=1
M685 550 563 559 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=120980 $D=1
M686 570 119 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=116350 $D=1
M687 571 559 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=120980 $D=1
M688 572 562 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=116350 $D=1
M689 573 563 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=120980 $D=1
M690 574 572 570 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=116350 $D=1
M691 575 573 571 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=120980 $D=1
M692 557 562 574 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=116350 $D=1
M693 558 563 575 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=120980 $D=1
M694 576 549 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=116350 $D=1
M695 577 550 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=120980 $D=1
M696 7 557 576 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=116350 $D=1
M697 8 558 577 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=120980 $D=1
M698 578 574 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=116350 $D=1
M699 579 575 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=120980 $D=1
M700 789 549 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=116350 $D=1
M701 790 550 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=120980 $D=1
M702 580 557 789 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=116350 $D=1
M703 581 558 790 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=120980 $D=1
M704 791 549 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=116350 $D=1
M705 792 550 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=120980 $D=1
M706 582 557 791 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=116350 $D=1
M707 583 558 792 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=120980 $D=1
M708 586 549 584 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=116350 $D=1
M709 587 550 585 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=120980 $D=1
M710 584 557 586 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=116350 $D=1
M711 585 558 587 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=120980 $D=1
M712 7 582 584 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=116350 $D=1
M713 8 583 585 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=120980 $D=1
M714 588 122 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=116350 $D=1
M715 589 122 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=120980 $D=1
M716 590 588 576 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=116350 $D=1
M717 591 589 577 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=120980 $D=1
M718 580 122 590 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=116350 $D=1
M719 581 122 591 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=120980 $D=1
M720 592 588 578 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=116350 $D=1
M721 593 589 579 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=120980 $D=1
M722 586 122 592 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=116350 $D=1
M723 587 122 593 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=120980 $D=1
M724 594 123 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=116350 $D=1
M725 595 123 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=120980 $D=1
M726 596 594 592 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=116350 $D=1
M727 597 595 593 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=120980 $D=1
M728 590 123 596 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=116350 $D=1
M729 591 123 597 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=120980 $D=1
M730 11 596 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=116350 $D=1
M731 12 597 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=120980 $D=1
M732 598 124 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=116350 $D=1
M733 599 124 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=120980 $D=1
M734 600 598 125 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=116350 $D=1
M735 601 599 126 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=120980 $D=1
M736 127 124 600 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=116350 $D=1
M737 128 124 601 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=120980 $D=1
M738 602 124 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=116350 $D=1
M739 603 124 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=120980 $D=1
M740 607 602 129 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=116350 $D=1
M741 608 603 131 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=120980 $D=1
M742 132 124 607 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=116350 $D=1
M743 130 124 608 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=120980 $D=1
M744 609 124 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=116350 $D=1
M745 610 124 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=120980 $D=1
M746 134 609 120 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=116350 $D=1
M747 134 610 133 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=120980 $D=1
M748 135 124 134 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=116350 $D=1
M749 136 124 134 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=120980 $D=1
M750 611 124 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=116350 $D=1
M751 612 124 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=120980 $D=1
M752 613 611 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=116350 $D=1
M753 614 612 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=120980 $D=1
M754 137 124 613 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=116350 $D=1
M755 138 124 614 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=120980 $D=1
M756 615 124 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=116350 $D=1
M757 616 124 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=120980 $D=1
M758 617 615 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=116350 $D=1
M759 618 616 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=120980 $D=1
M760 139 124 617 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=116350 $D=1
M761 140 124 618 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=120980 $D=1
M762 7 549 771 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=116350 $D=1
M763 8 550 772 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=120980 $D=1
M764 128 771 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=116350 $D=1
M765 125 772 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=120980 $D=1
M766 619 141 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=116350 $D=1
M767 620 141 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=120980 $D=1
M768 142 619 128 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=116350 $D=1
M769 143 620 125 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=120980 $D=1
M770 600 141 142 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=116350 $D=1
M771 601 141 143 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=120980 $D=1
M772 621 144 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=116350 $D=1
M773 622 144 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=120980 $D=1
M774 145 621 142 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=116350 $D=1
M775 146 622 143 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=120980 $D=1
M776 607 144 145 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=116350 $D=1
M777 608 144 146 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=120980 $D=1
M778 623 147 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=116350 $D=1
M779 624 147 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=120980 $D=1
M780 148 623 145 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=116350 $D=1
M781 149 624 146 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=120980 $D=1
M782 134 147 148 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=116350 $D=1
M783 134 147 149 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=120980 $D=1
M784 625 150 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=116350 $D=1
M785 626 150 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=120980 $D=1
M786 151 625 148 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=116350 $D=1
M787 152 626 149 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=120980 $D=1
M788 613 150 151 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=116350 $D=1
M789 614 150 152 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=120980 $D=1
M790 627 126 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=116350 $D=1
M791 628 126 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=120980 $D=1
M792 199 627 151 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=116350 $D=1
M793 200 628 152 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=120980 $D=1
M794 617 126 199 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=116350 $D=1
M795 618 126 200 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=120980 $D=1
M796 629 153 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=116350 $D=1
M797 630 153 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=120980 $D=1
M798 631 629 111 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=116350 $D=1
M799 632 630 112 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=120980 $D=1
M800 9 153 631 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=116350 $D=1
M801 10 153 632 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=120980 $D=1
M802 793 539 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=116350 $D=1
M803 794 540 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=120980 $D=1
M804 633 631 793 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=116350 $D=1
M805 634 632 794 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=120980 $D=1
M806 637 539 635 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=116350 $D=1
M807 638 540 636 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=120980 $D=1
M808 635 631 637 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=116350 $D=1
M809 636 632 638 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=120980 $D=1
M810 7 633 635 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=116350 $D=1
M811 8 634 636 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=120980 $D=1
M812 795 639 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=116350 $D=1
M813 796 640 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=120980 $D=1
M814 773 637 795 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=116350 $D=1
M815 774 638 796 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=120980 $D=1
M816 640 773 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=116350 $D=1
M817 154 774 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=120980 $D=1
M818 641 539 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=116350 $D=1
M819 642 540 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=120980 $D=1
M820 7 643 641 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=116350 $D=1
M821 8 644 642 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=120980 $D=1
M822 643 631 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=116350 $D=1
M823 644 632 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=120980 $D=1
M824 797 641 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=116350 $D=1
M825 798 642 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=120980 $D=1
M826 645 639 797 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=116350 $D=1
M827 646 640 798 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=120980 $D=1
M828 648 155 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=116350 $D=1
M829 649 647 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=120980 $D=1
M830 799 645 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=116350 $D=1
M831 800 646 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=120980 $D=1
M832 647 648 799 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=116350 $D=1
M833 156 649 800 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=120980 $D=1
M834 651 650 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=116350 $D=1
M835 652 157 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=120980 $D=1
M836 7 655 653 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=116350 $D=1
M837 8 656 654 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=120980 $D=1
M838 657 114 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=116350 $D=1
M839 658 115 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=120980 $D=1
M840 655 657 650 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=116350 $D=1
M841 656 658 157 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=120980 $D=1
M842 651 114 655 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=116350 $D=1
M843 652 115 656 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=120980 $D=1
M844 659 653 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=116350 $D=1
M845 660 654 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=120980 $D=1
M846 158 659 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=116350 $D=1
M847 650 660 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=120980 $D=1
M848 114 653 158 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=116350 $D=1
M849 115 654 650 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=120980 $D=1
M850 661 158 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=116350 $D=1
M851 662 650 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=120980 $D=1
M852 663 653 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=116350 $D=1
M853 664 654 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=120980 $D=1
M854 201 663 661 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=116350 $D=1
M855 202 664 662 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=120980 $D=1
M856 7 653 201 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=116350 $D=1
M857 8 654 202 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=120980 $D=1
M858 665 159 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=116350 $D=1
M859 666 159 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=120980 $D=1
M860 667 665 201 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=116350 $D=1
M861 668 666 202 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=120980 $D=1
M862 11 159 667 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=116350 $D=1
M863 12 159 668 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=120980 $D=1
M864 669 160 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=116350 $D=1
M865 670 160 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=120980 $D=1
M866 160 669 667 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=116350 $D=1
M867 160 670 668 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=120980 $D=1
M868 7 160 160 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=116350 $D=1
M869 8 160 160 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=120980 $D=1
M870 671 110 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=116350 $D=1
M871 672 110 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=120980 $D=1
M872 7 671 673 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=116350 $D=1
M873 8 672 674 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=120980 $D=1
M874 675 110 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=116350 $D=1
M875 676 110 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=120980 $D=1
M876 677 671 160 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=116350 $D=1
M877 678 672 160 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=120980 $D=1
M878 7 677 775 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=116350 $D=1
M879 8 678 776 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=120980 $D=1
M880 679 775 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=116350 $D=1
M881 680 776 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=120980 $D=1
M882 677 673 679 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=116350 $D=1
M883 678 674 680 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=120980 $D=1
M884 681 110 679 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=116350 $D=1
M885 682 110 680 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=120980 $D=1
M886 7 685 683 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=116350 $D=1
M887 8 686 684 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=120980 $D=1
M888 685 110 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=116350 $D=1
M889 686 110 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=120980 $D=1
M890 777 681 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=116350 $D=1
M891 778 682 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=120980 $D=1
M892 687 683 777 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=116350 $D=1
M893 688 684 778 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=120980 $D=1
M894 7 687 114 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=116350 $D=1
M895 8 688 115 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=120980 $D=1
M896 779 114 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=116350 $D=1
M897 780 115 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=120980 $D=1
M898 687 685 779 7 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=116350 $D=1
M899 688 686 780 8 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=120980 $D=1
M900 175 1 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=117600 $D=0
M901 176 1 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=122230 $D=0
M902 177 1 2 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=117600 $D=0
M903 178 1 3 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=122230 $D=0
M904 7 175 177 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=117600 $D=0
M905 8 176 178 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=122230 $D=0
M906 179 1 2 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=117600 $D=0
M907 180 1 3 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=122230 $D=0
M908 2 175 179 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=117600 $D=0
M909 3 176 180 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=122230 $D=0
M910 181 1 2 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=117600 $D=0
M911 182 1 3 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=122230 $D=0
M912 2 175 181 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=117600 $D=0
M913 3 176 182 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=122230 $D=0
M914 185 4 181 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=117600 $D=0
M915 186 4 182 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=122230 $D=0
M916 183 4 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=117600 $D=0
M917 184 4 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=122230 $D=0
M918 187 4 179 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=117600 $D=0
M919 188 4 180 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=122230 $D=0
M920 177 183 187 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=117600 $D=0
M921 178 184 188 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=122230 $D=0
M922 189 5 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=117600 $D=0
M923 190 5 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=122230 $D=0
M924 191 5 187 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=117600 $D=0
M925 192 5 188 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=122230 $D=0
M926 185 189 191 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=117600 $D=0
M927 186 190 192 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=122230 $D=0
M928 193 6 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=117600 $D=0
M929 194 6 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=122230 $D=0
M930 195 6 7 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=117600 $D=0
M931 196 6 8 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=122230 $D=0
M932 9 193 195 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=117600 $D=0
M933 10 194 196 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=122230 $D=0
M934 197 6 11 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=117600 $D=0
M935 198 6 12 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=122230 $D=0
M936 199 193 197 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=117600 $D=0
M937 200 194 198 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=122230 $D=0
M938 203 6 201 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=117600 $D=0
M939 204 6 202 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=122230 $D=0
M940 191 193 203 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=117600 $D=0
M941 192 194 204 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=122230 $D=0
M942 207 13 203 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=117600 $D=0
M943 208 13 204 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=122230 $D=0
M944 205 13 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=117600 $D=0
M945 206 13 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=122230 $D=0
M946 209 13 197 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=117600 $D=0
M947 210 13 198 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=122230 $D=0
M948 195 205 209 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=117600 $D=0
M949 196 206 210 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=122230 $D=0
M950 211 14 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=117600 $D=0
M951 212 14 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=122230 $D=0
M952 213 14 209 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=117600 $D=0
M953 214 14 210 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=122230 $D=0
M954 207 211 213 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=117600 $D=0
M955 208 212 214 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=122230 $D=0
M956 161 15 215 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=117600 $D=0
M957 162 15 216 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=122230 $D=0
M958 217 16 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=117600 $D=0
M959 218 16 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=122230 $D=0
M960 219 215 213 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=117600 $D=0
M961 220 216 214 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=122230 $D=0
M962 161 219 689 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=117600 $D=0
M963 162 220 690 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=122230 $D=0
M964 221 689 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=117600 $D=0
M965 222 690 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=122230 $D=0
M966 219 15 221 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=117600 $D=0
M967 220 15 222 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=122230 $D=0
M968 221 217 223 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=117600 $D=0
M969 222 218 224 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=122230 $D=0
M970 227 225 221 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=117600 $D=0
M971 228 226 222 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=122230 $D=0
M972 225 17 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=117600 $D=0
M973 226 17 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=122230 $D=0
M974 161 18 229 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=117600 $D=0
M975 162 18 230 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=122230 $D=0
M976 231 19 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=117600 $D=0
M977 232 19 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=122230 $D=0
M978 233 229 213 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=117600 $D=0
M979 234 230 214 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=122230 $D=0
M980 161 233 691 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=117600 $D=0
M981 162 234 692 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=122230 $D=0
M982 235 691 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=117600 $D=0
M983 236 692 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=122230 $D=0
M984 233 18 235 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=117600 $D=0
M985 234 18 236 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=122230 $D=0
M986 235 231 223 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=117600 $D=0
M987 236 232 224 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=122230 $D=0
M988 227 237 235 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=117600 $D=0
M989 228 238 236 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=122230 $D=0
M990 237 20 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=117600 $D=0
M991 238 20 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=122230 $D=0
M992 161 21 239 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=117600 $D=0
M993 162 21 240 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=122230 $D=0
M994 241 22 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=117600 $D=0
M995 242 22 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=122230 $D=0
M996 243 239 213 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=117600 $D=0
M997 244 240 214 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=122230 $D=0
M998 161 243 693 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=117600 $D=0
M999 162 244 694 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=122230 $D=0
M1000 245 693 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=117600 $D=0
M1001 246 694 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=122230 $D=0
M1002 243 21 245 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=117600 $D=0
M1003 244 21 246 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=122230 $D=0
M1004 245 241 223 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=117600 $D=0
M1005 246 242 224 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=122230 $D=0
M1006 227 247 245 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=117600 $D=0
M1007 228 248 246 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=122230 $D=0
M1008 247 23 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=117600 $D=0
M1009 248 23 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=122230 $D=0
M1010 161 24 249 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=117600 $D=0
M1011 162 24 250 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=122230 $D=0
M1012 251 25 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=117600 $D=0
M1013 252 25 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=122230 $D=0
M1014 253 249 213 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=117600 $D=0
M1015 254 250 214 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=122230 $D=0
M1016 161 253 695 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=117600 $D=0
M1017 162 254 696 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=122230 $D=0
M1018 255 695 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=117600 $D=0
M1019 256 696 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=122230 $D=0
M1020 253 24 255 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=117600 $D=0
M1021 254 24 256 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=122230 $D=0
M1022 255 251 223 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=117600 $D=0
M1023 256 252 224 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=122230 $D=0
M1024 227 257 255 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=117600 $D=0
M1025 228 258 256 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=122230 $D=0
M1026 257 26 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=117600 $D=0
M1027 258 26 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=122230 $D=0
M1028 161 27 259 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=117600 $D=0
M1029 162 27 260 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=122230 $D=0
M1030 261 28 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=117600 $D=0
M1031 262 28 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=122230 $D=0
M1032 263 259 213 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=117600 $D=0
M1033 264 260 214 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=122230 $D=0
M1034 161 263 697 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=117600 $D=0
M1035 162 264 698 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=122230 $D=0
M1036 265 697 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=117600 $D=0
M1037 266 698 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=122230 $D=0
M1038 263 27 265 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=117600 $D=0
M1039 264 27 266 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=122230 $D=0
M1040 265 261 223 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=117600 $D=0
M1041 266 262 224 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=122230 $D=0
M1042 227 267 265 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=117600 $D=0
M1043 228 268 266 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=122230 $D=0
M1044 267 29 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=117600 $D=0
M1045 268 29 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=122230 $D=0
M1046 161 30 269 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=117600 $D=0
M1047 162 30 270 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=122230 $D=0
M1048 271 31 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=117600 $D=0
M1049 272 31 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=122230 $D=0
M1050 273 269 213 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=117600 $D=0
M1051 274 270 214 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=122230 $D=0
M1052 161 273 699 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=117600 $D=0
M1053 162 274 700 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=122230 $D=0
M1054 275 699 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=117600 $D=0
M1055 276 700 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=122230 $D=0
M1056 273 30 275 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=117600 $D=0
M1057 274 30 276 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=122230 $D=0
M1058 275 271 223 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=117600 $D=0
M1059 276 272 224 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=122230 $D=0
M1060 227 277 275 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=117600 $D=0
M1061 228 278 276 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=122230 $D=0
M1062 277 32 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=117600 $D=0
M1063 278 32 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=122230 $D=0
M1064 161 33 279 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=117600 $D=0
M1065 162 33 280 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=122230 $D=0
M1066 281 34 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=117600 $D=0
M1067 282 34 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=122230 $D=0
M1068 283 279 213 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=117600 $D=0
M1069 284 280 214 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=122230 $D=0
M1070 161 283 701 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=117600 $D=0
M1071 162 284 702 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=122230 $D=0
M1072 285 701 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=117600 $D=0
M1073 286 702 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=122230 $D=0
M1074 283 33 285 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=117600 $D=0
M1075 284 33 286 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=122230 $D=0
M1076 285 281 223 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=117600 $D=0
M1077 286 282 224 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=122230 $D=0
M1078 227 287 285 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=117600 $D=0
M1079 228 288 286 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=122230 $D=0
M1080 287 35 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=117600 $D=0
M1081 288 35 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=122230 $D=0
M1082 161 36 289 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=117600 $D=0
M1083 162 36 290 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=122230 $D=0
M1084 291 37 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=117600 $D=0
M1085 292 37 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=122230 $D=0
M1086 293 289 213 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=117600 $D=0
M1087 294 290 214 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=122230 $D=0
M1088 161 293 703 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=117600 $D=0
M1089 162 294 704 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=122230 $D=0
M1090 295 703 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=117600 $D=0
M1091 296 704 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=122230 $D=0
M1092 293 36 295 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=117600 $D=0
M1093 294 36 296 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=122230 $D=0
M1094 295 291 223 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=117600 $D=0
M1095 296 292 224 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=122230 $D=0
M1096 227 297 295 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=117600 $D=0
M1097 228 298 296 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=122230 $D=0
M1098 297 38 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=117600 $D=0
M1099 298 38 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=122230 $D=0
M1100 161 39 299 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=117600 $D=0
M1101 162 39 300 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=122230 $D=0
M1102 301 40 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=117600 $D=0
M1103 302 40 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=122230 $D=0
M1104 303 299 213 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=117600 $D=0
M1105 304 300 214 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=122230 $D=0
M1106 161 303 705 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=117600 $D=0
M1107 162 304 706 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=122230 $D=0
M1108 305 705 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=117600 $D=0
M1109 306 706 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=122230 $D=0
M1110 303 39 305 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=117600 $D=0
M1111 304 39 306 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=122230 $D=0
M1112 305 301 223 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=117600 $D=0
M1113 306 302 224 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=122230 $D=0
M1114 227 307 305 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=117600 $D=0
M1115 228 308 306 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=122230 $D=0
M1116 307 41 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=117600 $D=0
M1117 308 41 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=122230 $D=0
M1118 161 42 309 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=117600 $D=0
M1119 162 42 310 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=122230 $D=0
M1120 311 43 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=117600 $D=0
M1121 312 43 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=122230 $D=0
M1122 313 309 213 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=117600 $D=0
M1123 314 310 214 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=122230 $D=0
M1124 161 313 707 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=117600 $D=0
M1125 162 314 708 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=122230 $D=0
M1126 315 707 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=117600 $D=0
M1127 316 708 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=122230 $D=0
M1128 313 42 315 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=117600 $D=0
M1129 314 42 316 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=122230 $D=0
M1130 315 311 223 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=117600 $D=0
M1131 316 312 224 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=122230 $D=0
M1132 227 317 315 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=117600 $D=0
M1133 228 318 316 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=122230 $D=0
M1134 317 44 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=117600 $D=0
M1135 318 44 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=122230 $D=0
M1136 161 45 319 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=117600 $D=0
M1137 162 45 320 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=122230 $D=0
M1138 321 46 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=117600 $D=0
M1139 322 46 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=122230 $D=0
M1140 323 319 213 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=117600 $D=0
M1141 324 320 214 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=122230 $D=0
M1142 161 323 709 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=117600 $D=0
M1143 162 324 710 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=122230 $D=0
M1144 325 709 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=117600 $D=0
M1145 326 710 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=122230 $D=0
M1146 323 45 325 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=117600 $D=0
M1147 324 45 326 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=122230 $D=0
M1148 325 321 223 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=117600 $D=0
M1149 326 322 224 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=122230 $D=0
M1150 227 327 325 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=117600 $D=0
M1151 228 328 326 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=122230 $D=0
M1152 327 47 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=117600 $D=0
M1153 328 47 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=122230 $D=0
M1154 161 48 329 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=117600 $D=0
M1155 162 48 330 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=122230 $D=0
M1156 331 49 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=117600 $D=0
M1157 332 49 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=122230 $D=0
M1158 333 329 213 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=117600 $D=0
M1159 334 330 214 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=122230 $D=0
M1160 161 333 711 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=117600 $D=0
M1161 162 334 712 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=122230 $D=0
M1162 335 711 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=117600 $D=0
M1163 336 712 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=122230 $D=0
M1164 333 48 335 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=117600 $D=0
M1165 334 48 336 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=122230 $D=0
M1166 335 331 223 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=117600 $D=0
M1167 336 332 224 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=122230 $D=0
M1168 227 337 335 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=117600 $D=0
M1169 228 338 336 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=122230 $D=0
M1170 337 50 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=117600 $D=0
M1171 338 50 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=122230 $D=0
M1172 161 51 339 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=117600 $D=0
M1173 162 51 340 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=122230 $D=0
M1174 341 52 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=117600 $D=0
M1175 342 52 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=122230 $D=0
M1176 343 339 213 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=117600 $D=0
M1177 344 340 214 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=122230 $D=0
M1178 161 343 713 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=117600 $D=0
M1179 162 344 714 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=122230 $D=0
M1180 345 713 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=117600 $D=0
M1181 346 714 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=122230 $D=0
M1182 343 51 345 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=117600 $D=0
M1183 344 51 346 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=122230 $D=0
M1184 345 341 223 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=117600 $D=0
M1185 346 342 224 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=122230 $D=0
M1186 227 347 345 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=117600 $D=0
M1187 228 348 346 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=122230 $D=0
M1188 347 53 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=117600 $D=0
M1189 348 53 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=122230 $D=0
M1190 161 54 349 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=117600 $D=0
M1191 162 54 350 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=122230 $D=0
M1192 351 55 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=117600 $D=0
M1193 352 55 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=122230 $D=0
M1194 353 349 213 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=117600 $D=0
M1195 354 350 214 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=122230 $D=0
M1196 161 353 715 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=117600 $D=0
M1197 162 354 716 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=122230 $D=0
M1198 355 715 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=117600 $D=0
M1199 356 716 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=122230 $D=0
M1200 353 54 355 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=117600 $D=0
M1201 354 54 356 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=122230 $D=0
M1202 355 351 223 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=117600 $D=0
M1203 356 352 224 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=122230 $D=0
M1204 227 357 355 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=117600 $D=0
M1205 228 358 356 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=122230 $D=0
M1206 357 56 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=117600 $D=0
M1207 358 56 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=122230 $D=0
M1208 161 57 359 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=117600 $D=0
M1209 162 57 360 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=122230 $D=0
M1210 361 58 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=117600 $D=0
M1211 362 58 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=122230 $D=0
M1212 363 359 213 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=117600 $D=0
M1213 364 360 214 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=122230 $D=0
M1214 161 363 717 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=117600 $D=0
M1215 162 364 718 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=122230 $D=0
M1216 365 717 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=117600 $D=0
M1217 366 718 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=122230 $D=0
M1218 363 57 365 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=117600 $D=0
M1219 364 57 366 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=122230 $D=0
M1220 365 361 223 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=117600 $D=0
M1221 366 362 224 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=122230 $D=0
M1222 227 367 365 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=117600 $D=0
M1223 228 368 366 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=122230 $D=0
M1224 367 59 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=117600 $D=0
M1225 368 59 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=122230 $D=0
M1226 161 60 369 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=117600 $D=0
M1227 162 60 370 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=122230 $D=0
M1228 371 61 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=117600 $D=0
M1229 372 61 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=122230 $D=0
M1230 373 369 213 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=117600 $D=0
M1231 374 370 214 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=122230 $D=0
M1232 161 373 719 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=117600 $D=0
M1233 162 374 720 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=122230 $D=0
M1234 375 719 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=117600 $D=0
M1235 376 720 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=122230 $D=0
M1236 373 60 375 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=117600 $D=0
M1237 374 60 376 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=122230 $D=0
M1238 375 371 223 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=117600 $D=0
M1239 376 372 224 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=122230 $D=0
M1240 227 377 375 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=117600 $D=0
M1241 228 378 376 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=122230 $D=0
M1242 377 62 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=117600 $D=0
M1243 378 62 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=122230 $D=0
M1244 161 63 379 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=117600 $D=0
M1245 162 63 380 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=122230 $D=0
M1246 381 64 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=117600 $D=0
M1247 382 64 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=122230 $D=0
M1248 383 379 213 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=117600 $D=0
M1249 384 380 214 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=122230 $D=0
M1250 161 383 721 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=117600 $D=0
M1251 162 384 722 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=122230 $D=0
M1252 385 721 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=117600 $D=0
M1253 386 722 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=122230 $D=0
M1254 383 63 385 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=117600 $D=0
M1255 384 63 386 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=122230 $D=0
M1256 385 381 223 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=117600 $D=0
M1257 386 382 224 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=122230 $D=0
M1258 227 387 385 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=117600 $D=0
M1259 228 388 386 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=122230 $D=0
M1260 387 65 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=117600 $D=0
M1261 388 65 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=122230 $D=0
M1262 161 66 389 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=117600 $D=0
M1263 162 66 390 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=122230 $D=0
M1264 391 67 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=117600 $D=0
M1265 392 67 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=122230 $D=0
M1266 393 389 213 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=117600 $D=0
M1267 394 390 214 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=122230 $D=0
M1268 161 393 723 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=117600 $D=0
M1269 162 394 724 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=122230 $D=0
M1270 395 723 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=117600 $D=0
M1271 396 724 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=122230 $D=0
M1272 393 66 395 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=117600 $D=0
M1273 394 66 396 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=122230 $D=0
M1274 395 391 223 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=117600 $D=0
M1275 396 392 224 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=122230 $D=0
M1276 227 397 395 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=117600 $D=0
M1277 228 398 396 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=122230 $D=0
M1278 397 68 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=117600 $D=0
M1279 398 68 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=122230 $D=0
M1280 161 69 399 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=117600 $D=0
M1281 162 69 400 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=122230 $D=0
M1282 401 70 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=117600 $D=0
M1283 402 70 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=122230 $D=0
M1284 403 399 213 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=117600 $D=0
M1285 404 400 214 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=122230 $D=0
M1286 161 403 725 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=117600 $D=0
M1287 162 404 726 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=122230 $D=0
M1288 405 725 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=117600 $D=0
M1289 406 726 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=122230 $D=0
M1290 403 69 405 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=117600 $D=0
M1291 404 69 406 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=122230 $D=0
M1292 405 401 223 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=117600 $D=0
M1293 406 402 224 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=122230 $D=0
M1294 227 407 405 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=117600 $D=0
M1295 228 408 406 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=122230 $D=0
M1296 407 71 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=117600 $D=0
M1297 408 71 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=122230 $D=0
M1298 161 72 409 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=117600 $D=0
M1299 162 72 410 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=122230 $D=0
M1300 411 73 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=117600 $D=0
M1301 412 73 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=122230 $D=0
M1302 413 409 213 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=117600 $D=0
M1303 414 410 214 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=122230 $D=0
M1304 161 413 727 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=117600 $D=0
M1305 162 414 728 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=122230 $D=0
M1306 415 727 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=117600 $D=0
M1307 416 728 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=122230 $D=0
M1308 413 72 415 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=117600 $D=0
M1309 414 72 416 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=122230 $D=0
M1310 415 411 223 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=117600 $D=0
M1311 416 412 224 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=122230 $D=0
M1312 227 417 415 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=117600 $D=0
M1313 228 418 416 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=122230 $D=0
M1314 417 74 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=117600 $D=0
M1315 418 74 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=122230 $D=0
M1316 161 75 419 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=117600 $D=0
M1317 162 75 420 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=122230 $D=0
M1318 421 76 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=117600 $D=0
M1319 422 76 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=122230 $D=0
M1320 423 419 213 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=117600 $D=0
M1321 424 420 214 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=122230 $D=0
M1322 161 423 729 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=117600 $D=0
M1323 162 424 730 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=122230 $D=0
M1324 425 729 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=117600 $D=0
M1325 426 730 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=122230 $D=0
M1326 423 75 425 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=117600 $D=0
M1327 424 75 426 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=122230 $D=0
M1328 425 421 223 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=117600 $D=0
M1329 426 422 224 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=122230 $D=0
M1330 227 427 425 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=117600 $D=0
M1331 228 428 426 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=122230 $D=0
M1332 427 77 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=117600 $D=0
M1333 428 77 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=122230 $D=0
M1334 161 78 429 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=117600 $D=0
M1335 162 78 430 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=122230 $D=0
M1336 431 79 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=117600 $D=0
M1337 432 79 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=122230 $D=0
M1338 433 429 213 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=117600 $D=0
M1339 434 430 214 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=122230 $D=0
M1340 161 433 731 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=117600 $D=0
M1341 162 434 732 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=122230 $D=0
M1342 435 731 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=117600 $D=0
M1343 436 732 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=122230 $D=0
M1344 433 78 435 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=117600 $D=0
M1345 434 78 436 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=122230 $D=0
M1346 435 431 223 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=117600 $D=0
M1347 436 432 224 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=122230 $D=0
M1348 227 437 435 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=117600 $D=0
M1349 228 438 436 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=122230 $D=0
M1350 437 80 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=117600 $D=0
M1351 438 80 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=122230 $D=0
M1352 161 81 439 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=117600 $D=0
M1353 162 81 440 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=122230 $D=0
M1354 441 82 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=117600 $D=0
M1355 442 82 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=122230 $D=0
M1356 443 439 213 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=117600 $D=0
M1357 444 440 214 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=122230 $D=0
M1358 161 443 733 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=117600 $D=0
M1359 162 444 734 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=122230 $D=0
M1360 445 733 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=117600 $D=0
M1361 446 734 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=122230 $D=0
M1362 443 81 445 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=117600 $D=0
M1363 444 81 446 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=122230 $D=0
M1364 445 441 223 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=117600 $D=0
M1365 446 442 224 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=122230 $D=0
M1366 227 447 445 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=117600 $D=0
M1367 228 448 446 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=122230 $D=0
M1368 447 83 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=117600 $D=0
M1369 448 83 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=122230 $D=0
M1370 161 84 449 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=117600 $D=0
M1371 162 84 450 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=122230 $D=0
M1372 451 85 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=117600 $D=0
M1373 452 85 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=122230 $D=0
M1374 453 449 213 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=117600 $D=0
M1375 454 450 214 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=122230 $D=0
M1376 161 453 735 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=117600 $D=0
M1377 162 454 736 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=122230 $D=0
M1378 455 735 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=117600 $D=0
M1379 456 736 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=122230 $D=0
M1380 453 84 455 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=117600 $D=0
M1381 454 84 456 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=122230 $D=0
M1382 455 451 223 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=117600 $D=0
M1383 456 452 224 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=122230 $D=0
M1384 227 457 455 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=117600 $D=0
M1385 228 458 456 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=122230 $D=0
M1386 457 86 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=117600 $D=0
M1387 458 86 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=122230 $D=0
M1388 161 87 459 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=117600 $D=0
M1389 162 87 460 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=122230 $D=0
M1390 461 88 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=117600 $D=0
M1391 462 88 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=122230 $D=0
M1392 463 459 213 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=117600 $D=0
M1393 464 460 214 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=122230 $D=0
M1394 161 463 737 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=117600 $D=0
M1395 162 464 738 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=122230 $D=0
M1396 465 737 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=117600 $D=0
M1397 466 738 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=122230 $D=0
M1398 463 87 465 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=117600 $D=0
M1399 464 87 466 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=122230 $D=0
M1400 465 461 223 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=117600 $D=0
M1401 466 462 224 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=122230 $D=0
M1402 227 467 465 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=117600 $D=0
M1403 228 468 466 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=122230 $D=0
M1404 467 89 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=117600 $D=0
M1405 468 89 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=122230 $D=0
M1406 161 90 469 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=117600 $D=0
M1407 162 90 470 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=122230 $D=0
M1408 471 91 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=117600 $D=0
M1409 472 91 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=122230 $D=0
M1410 473 469 213 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=117600 $D=0
M1411 474 470 214 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=122230 $D=0
M1412 161 473 739 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=117600 $D=0
M1413 162 474 740 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=122230 $D=0
M1414 475 739 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=117600 $D=0
M1415 476 740 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=122230 $D=0
M1416 473 90 475 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=117600 $D=0
M1417 474 90 476 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=122230 $D=0
M1418 475 471 223 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=117600 $D=0
M1419 476 472 224 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=122230 $D=0
M1420 227 477 475 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=117600 $D=0
M1421 228 478 476 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=122230 $D=0
M1422 477 92 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=117600 $D=0
M1423 478 92 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=122230 $D=0
M1424 161 93 479 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=117600 $D=0
M1425 162 93 480 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=122230 $D=0
M1426 481 94 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=117600 $D=0
M1427 482 94 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=122230 $D=0
M1428 483 479 213 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=117600 $D=0
M1429 484 480 214 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=122230 $D=0
M1430 161 483 741 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=117600 $D=0
M1431 162 484 742 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=122230 $D=0
M1432 485 741 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=117600 $D=0
M1433 486 742 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=122230 $D=0
M1434 483 93 485 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=117600 $D=0
M1435 484 93 486 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=122230 $D=0
M1436 485 481 223 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=117600 $D=0
M1437 486 482 224 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=122230 $D=0
M1438 227 487 485 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=117600 $D=0
M1439 228 488 486 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=122230 $D=0
M1440 487 95 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=117600 $D=0
M1441 488 95 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=122230 $D=0
M1442 161 96 489 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=117600 $D=0
M1443 162 96 490 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=122230 $D=0
M1444 491 97 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=117600 $D=0
M1445 492 97 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=122230 $D=0
M1446 493 489 213 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=117600 $D=0
M1447 494 490 214 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=122230 $D=0
M1448 161 493 743 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=117600 $D=0
M1449 162 494 744 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=122230 $D=0
M1450 495 743 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=117600 $D=0
M1451 496 744 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=122230 $D=0
M1452 493 96 495 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=117600 $D=0
M1453 494 96 496 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=122230 $D=0
M1454 495 491 223 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=117600 $D=0
M1455 496 492 224 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=122230 $D=0
M1456 227 497 495 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=117600 $D=0
M1457 228 498 496 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=122230 $D=0
M1458 497 98 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=117600 $D=0
M1459 498 98 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=122230 $D=0
M1460 161 99 499 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=117600 $D=0
M1461 162 99 500 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=122230 $D=0
M1462 501 100 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=117600 $D=0
M1463 502 100 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=122230 $D=0
M1464 503 499 213 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=117600 $D=0
M1465 504 500 214 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=122230 $D=0
M1466 161 503 745 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=117600 $D=0
M1467 162 504 746 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=122230 $D=0
M1468 505 745 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=117600 $D=0
M1469 506 746 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=122230 $D=0
M1470 503 99 505 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=117600 $D=0
M1471 504 99 506 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=122230 $D=0
M1472 505 501 223 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=117600 $D=0
M1473 506 502 224 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=122230 $D=0
M1474 227 507 505 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=117600 $D=0
M1475 228 508 506 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=122230 $D=0
M1476 507 101 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=117600 $D=0
M1477 508 101 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=122230 $D=0
M1478 161 102 509 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=117600 $D=0
M1479 162 102 510 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=122230 $D=0
M1480 511 103 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=117600 $D=0
M1481 512 103 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=122230 $D=0
M1482 513 509 213 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=117600 $D=0
M1483 514 510 214 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=122230 $D=0
M1484 161 513 747 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=117600 $D=0
M1485 162 514 748 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=122230 $D=0
M1486 515 747 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=117600 $D=0
M1487 516 748 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=122230 $D=0
M1488 513 102 515 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=117600 $D=0
M1489 514 102 516 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=122230 $D=0
M1490 515 511 223 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=117600 $D=0
M1491 516 512 224 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=122230 $D=0
M1492 227 517 515 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=117600 $D=0
M1493 228 518 516 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=122230 $D=0
M1494 517 104 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=117600 $D=0
M1495 518 104 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=122230 $D=0
M1496 161 105 519 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=117600 $D=0
M1497 162 105 520 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=122230 $D=0
M1498 521 106 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=117600 $D=0
M1499 522 106 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=122230 $D=0
M1500 523 519 213 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=117600 $D=0
M1501 524 520 214 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=122230 $D=0
M1502 161 523 749 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=117600 $D=0
M1503 162 524 750 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=122230 $D=0
M1504 525 749 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=117600 $D=0
M1505 526 750 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=122230 $D=0
M1506 523 105 525 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=117600 $D=0
M1507 524 105 526 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=122230 $D=0
M1508 525 521 223 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=117600 $D=0
M1509 526 522 224 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=122230 $D=0
M1510 227 527 525 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=117600 $D=0
M1511 228 528 526 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=122230 $D=0
M1512 527 107 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=117600 $D=0
M1513 528 107 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=122230 $D=0
M1514 161 108 529 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=117600 $D=0
M1515 162 108 530 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=122230 $D=0
M1516 531 109 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=117600 $D=0
M1517 532 109 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=122230 $D=0
M1518 7 531 223 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=117600 $D=0
M1519 8 532 224 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=122230 $D=0
M1520 227 529 7 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=117600 $D=0
M1521 228 530 8 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=122230 $D=0
M1522 161 535 533 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=117600 $D=0
M1523 162 536 534 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=122230 $D=0
M1524 535 110 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=117600 $D=0
M1525 536 110 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=122230 $D=0
M1526 751 223 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=117600 $D=0
M1527 752 224 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=122230 $D=0
M1528 537 535 751 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=117600 $D=0
M1529 538 536 752 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=122230 $D=0
M1530 161 537 539 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=117600 $D=0
M1531 162 538 540 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=122230 $D=0
M1532 753 539 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=117600 $D=0
M1533 754 540 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=122230 $D=0
M1534 537 533 753 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=117600 $D=0
M1535 538 534 754 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=122230 $D=0
M1536 161 543 541 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=117600 $D=0
M1537 162 544 542 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=122230 $D=0
M1538 543 110 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=117600 $D=0
M1539 544 110 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=122230 $D=0
M1540 755 227 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=117600 $D=0
M1541 756 228 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=122230 $D=0
M1542 545 543 755 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=117600 $D=0
M1543 546 544 756 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=122230 $D=0
M1544 161 545 111 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=117600 $D=0
M1545 162 546 112 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=122230 $D=0
M1546 757 111 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=117600 $D=0
M1547 758 112 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=122230 $D=0
M1548 545 541 757 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=117600 $D=0
M1549 546 542 758 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=122230 $D=0
M1550 547 113 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=117600 $D=0
M1551 548 113 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=122230 $D=0
M1552 549 113 539 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=117600 $D=0
M1553 550 113 540 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=122230 $D=0
M1554 114 547 549 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=117600 $D=0
M1555 115 548 550 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=122230 $D=0
M1556 551 116 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=117600 $D=0
M1557 552 116 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=122230 $D=0
M1558 553 116 111 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=117600 $D=0
M1559 554 116 112 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=122230 $D=0
M1560 759 551 553 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=117600 $D=0
M1561 760 552 554 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=122230 $D=0
M1562 161 111 759 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=117600 $D=0
M1563 162 112 760 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=122230 $D=0
M1564 555 117 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=117600 $D=0
M1565 556 117 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=122230 $D=0
M1566 557 117 553 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=117600 $D=0
M1567 558 117 554 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=122230 $D=0
M1568 9 555 557 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=117600 $D=0
M1569 10 556 558 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=122230 $D=0
M1570 560 559 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=117600 $D=0
M1571 561 118 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=122230 $D=0
M1572 161 564 562 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=117600 $D=0
M1573 162 565 563 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=122230 $D=0
M1574 566 549 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=117600 $D=0
M1575 567 550 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=122230 $D=0
M1576 564 549 559 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=117600 $D=0
M1577 565 550 118 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=122230 $D=0
M1578 560 566 564 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=117600 $D=0
M1579 561 567 565 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=122230 $D=0
M1580 568 562 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=117600 $D=0
M1581 569 563 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=122230 $D=0
M1582 119 562 557 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=117600 $D=0
M1583 559 563 558 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=122230 $D=0
M1584 549 568 119 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=117600 $D=0
M1585 550 569 559 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=122230 $D=0
M1586 570 119 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=117600 $D=0
M1587 571 559 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=122230 $D=0
M1588 572 562 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=117600 $D=0
M1589 573 563 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=122230 $D=0
M1590 574 562 570 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=117600 $D=0
M1591 575 563 571 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=122230 $D=0
M1592 557 572 574 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=117600 $D=0
M1593 558 573 575 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=122230 $D=0
M1594 781 549 161 161 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=117240 $D=0
M1595 782 550 162 162 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=121870 $D=0
M1596 576 557 781 161 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=117240 $D=0
M1597 577 558 782 162 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=121870 $D=0
M1598 578 574 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=117600 $D=0
M1599 579 575 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=122230 $D=0
M1600 580 549 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=117600 $D=0
M1601 581 550 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=122230 $D=0
M1602 161 557 580 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=117600 $D=0
M1603 162 558 581 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=122230 $D=0
M1604 582 549 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=117600 $D=0
M1605 583 550 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=122230 $D=0
M1606 161 557 582 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=117600 $D=0
M1607 162 558 583 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=122230 $D=0
M1608 783 549 161 161 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=117420 $D=0
M1609 784 550 162 162 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=122050 $D=0
M1610 586 557 783 161 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=117420 $D=0
M1611 587 558 784 162 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=122050 $D=0
M1612 161 582 586 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=117600 $D=0
M1613 162 583 587 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=122230 $D=0
M1614 588 122 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=117600 $D=0
M1615 589 122 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=122230 $D=0
M1616 590 122 576 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=117600 $D=0
M1617 591 122 577 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=122230 $D=0
M1618 580 588 590 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=117600 $D=0
M1619 581 589 591 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=122230 $D=0
M1620 592 122 578 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=117600 $D=0
M1621 593 122 579 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=122230 $D=0
M1622 586 588 592 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=117600 $D=0
M1623 587 589 593 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=122230 $D=0
M1624 594 123 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=117600 $D=0
M1625 595 123 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=122230 $D=0
M1626 596 123 592 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=117600 $D=0
M1627 597 123 593 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=122230 $D=0
M1628 590 594 596 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=117600 $D=0
M1629 591 595 597 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=122230 $D=0
M1630 11 596 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=117600 $D=0
M1631 12 597 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=122230 $D=0
M1632 598 124 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=117600 $D=0
M1633 599 124 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=122230 $D=0
M1634 600 124 125 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=117600 $D=0
M1635 601 124 126 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=122230 $D=0
M1636 127 598 600 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=117600 $D=0
M1637 128 599 601 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=122230 $D=0
M1638 602 124 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=117600 $D=0
M1639 603 124 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=122230 $D=0
M1640 607 124 129 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=117600 $D=0
M1641 608 124 131 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=122230 $D=0
M1642 132 602 607 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=117600 $D=0
M1643 130 603 608 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=122230 $D=0
M1644 609 124 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=117600 $D=0
M1645 610 124 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=122230 $D=0
M1646 134 124 120 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=117600 $D=0
M1647 134 124 133 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=122230 $D=0
M1648 135 609 134 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=117600 $D=0
M1649 136 610 134 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=122230 $D=0
M1650 611 124 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=117600 $D=0
M1651 612 124 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=122230 $D=0
M1652 613 124 7 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=117600 $D=0
M1653 614 124 8 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=122230 $D=0
M1654 137 611 613 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=117600 $D=0
M1655 138 612 614 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=122230 $D=0
M1656 615 124 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=117600 $D=0
M1657 616 124 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=122230 $D=0
M1658 617 124 7 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=117600 $D=0
M1659 618 124 8 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=122230 $D=0
M1660 139 615 617 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=117600 $D=0
M1661 140 616 618 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=122230 $D=0
M1662 161 549 771 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=117600 $D=0
M1663 162 550 772 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=122230 $D=0
M1664 128 771 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=117600 $D=0
M1665 125 772 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=122230 $D=0
M1666 619 141 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=117600 $D=0
M1667 620 141 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=122230 $D=0
M1668 142 141 128 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=117600 $D=0
M1669 143 141 125 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=122230 $D=0
M1670 600 619 142 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=117600 $D=0
M1671 601 620 143 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=122230 $D=0
M1672 621 144 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=117600 $D=0
M1673 622 144 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=122230 $D=0
M1674 145 144 142 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=117600 $D=0
M1675 146 144 143 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=122230 $D=0
M1676 607 621 145 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=117600 $D=0
M1677 608 622 146 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=122230 $D=0
M1678 623 147 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=117600 $D=0
M1679 624 147 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=122230 $D=0
M1680 148 147 145 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=117600 $D=0
M1681 149 147 146 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=122230 $D=0
M1682 134 623 148 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=117600 $D=0
M1683 134 624 149 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=122230 $D=0
M1684 625 150 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=117600 $D=0
M1685 626 150 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=122230 $D=0
M1686 151 150 148 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=117600 $D=0
M1687 152 150 149 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=122230 $D=0
M1688 613 625 151 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=117600 $D=0
M1689 614 626 152 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=122230 $D=0
M1690 627 126 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=117600 $D=0
M1691 628 126 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=122230 $D=0
M1692 199 126 151 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=117600 $D=0
M1693 200 126 152 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=122230 $D=0
M1694 617 627 199 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=117600 $D=0
M1695 618 628 200 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=122230 $D=0
M1696 629 153 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=117600 $D=0
M1697 630 153 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=122230 $D=0
M1698 631 153 111 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=117600 $D=0
M1699 632 153 112 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=122230 $D=0
M1700 9 629 631 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=117600 $D=0
M1701 10 630 632 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=122230 $D=0
M1702 633 539 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=117600 $D=0
M1703 634 540 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=122230 $D=0
M1704 161 631 633 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=117600 $D=0
M1705 162 632 634 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=122230 $D=0
M1706 785 539 161 161 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=117420 $D=0
M1707 786 540 162 162 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=122050 $D=0
M1708 637 631 785 161 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=117420 $D=0
M1709 638 632 786 162 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=122050 $D=0
M1710 161 633 637 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=117600 $D=0
M1711 162 634 638 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=122230 $D=0
M1712 773 639 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=117600 $D=0
M1713 774 640 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=122230 $D=0
M1714 161 637 773 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=117600 $D=0
M1715 162 638 774 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=122230 $D=0
M1716 640 773 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=117600 $D=0
M1717 154 774 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=122230 $D=0
M1718 787 539 161 161 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=117240 $D=0
M1719 788 540 162 162 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=121870 $D=0
M1720 641 643 787 161 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=117240 $D=0
M1721 642 644 788 162 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=121870 $D=0
M1722 643 631 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=117600 $D=0
M1723 644 632 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=122230 $D=0
M1724 645 641 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=117600 $D=0
M1725 646 642 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=122230 $D=0
M1726 161 639 645 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=117600 $D=0
M1727 162 640 646 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=122230 $D=0
M1728 648 155 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=117600 $D=0
M1729 649 647 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=122230 $D=0
M1730 647 645 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=117600 $D=0
M1731 156 646 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=122230 $D=0
M1732 161 648 647 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=117600 $D=0
M1733 162 649 156 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=122230 $D=0
M1734 651 650 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=117600 $D=0
M1735 652 157 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=122230 $D=0
M1736 161 655 653 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=117600 $D=0
M1737 162 656 654 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=122230 $D=0
M1738 657 114 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=117600 $D=0
M1739 658 115 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=122230 $D=0
M1740 655 114 650 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=117600 $D=0
M1741 656 115 157 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=122230 $D=0
M1742 651 657 655 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=117600 $D=0
M1743 652 658 656 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=122230 $D=0
M1744 659 653 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=117600 $D=0
M1745 660 654 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=122230 $D=0
M1746 158 653 7 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=117600 $D=0
M1747 650 654 8 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=122230 $D=0
M1748 114 659 158 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=117600 $D=0
M1749 115 660 650 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=122230 $D=0
M1750 661 158 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=117600 $D=0
M1751 662 650 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=122230 $D=0
M1752 663 653 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=117600 $D=0
M1753 664 654 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=122230 $D=0
M1754 201 653 661 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=117600 $D=0
M1755 202 654 662 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=122230 $D=0
M1756 7 663 201 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=117600 $D=0
M1757 8 664 202 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=122230 $D=0
M1758 665 159 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=117600 $D=0
M1759 666 159 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=122230 $D=0
M1760 667 159 201 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=117600 $D=0
M1761 668 159 202 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=122230 $D=0
M1762 11 665 667 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=117600 $D=0
M1763 12 666 668 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=122230 $D=0
M1764 669 160 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=117600 $D=0
M1765 670 160 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=122230 $D=0
M1766 160 160 667 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=117600 $D=0
M1767 160 160 668 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=122230 $D=0
M1768 7 669 160 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=117600 $D=0
M1769 8 670 160 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=122230 $D=0
M1770 671 110 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=117600 $D=0
M1771 672 110 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=122230 $D=0
M1772 161 671 673 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=117600 $D=0
M1773 162 672 674 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=122230 $D=0
M1774 675 110 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=117600 $D=0
M1775 676 110 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=122230 $D=0
M1776 677 673 160 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=117600 $D=0
M1777 678 674 160 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=122230 $D=0
M1778 161 677 775 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=117600 $D=0
M1779 162 678 776 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=122230 $D=0
M1780 679 775 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=117600 $D=0
M1781 680 776 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=122230 $D=0
M1782 677 671 679 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=117600 $D=0
M1783 678 672 680 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=122230 $D=0
M1784 681 675 679 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=117600 $D=0
M1785 682 676 680 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=122230 $D=0
M1786 161 685 683 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=117600 $D=0
M1787 162 686 684 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=122230 $D=0
M1788 685 110 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=117600 $D=0
M1789 686 110 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=122230 $D=0
M1790 777 681 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=117600 $D=0
M1791 778 682 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=122230 $D=0
M1792 687 685 777 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=117600 $D=0
M1793 688 686 778 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=122230 $D=0
M1794 161 687 114 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=117600 $D=0
M1795 162 688 115 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=122230 $D=0
M1796 779 114 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=117600 $D=0
M1797 780 115 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=122230 $D=0
M1798 687 683 779 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=117600 $D=0
M1799 688 684 780 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=122230 $D=0
.ENDS
***************************************
.SUBCKT ICV_27 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162
** N=807 EP=162 IP=1514 FDC=1800
M0 179 1 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=107090 $D=1
M1 180 1 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=111720 $D=1
M2 181 179 2 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=107090 $D=1
M3 182 180 3 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=111720 $D=1
M4 4 1 181 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=107090 $D=1
M5 8 1 182 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=111720 $D=1
M6 183 179 3 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=107090 $D=1
M7 184 180 3 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=111720 $D=1
M8 2 1 183 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=107090 $D=1
M9 3 1 184 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=111720 $D=1
M10 185 179 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=107090 $D=1
M11 186 180 3 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=111720 $D=1
M12 2 1 185 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=107090 $D=1
M13 3 1 186 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=111720 $D=1
M14 189 187 185 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=107090 $D=1
M15 190 188 186 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=111720 $D=1
M16 187 5 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=107090 $D=1
M17 188 5 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=111720 $D=1
M18 191 187 183 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=107090 $D=1
M19 192 188 184 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=111720 $D=1
M20 181 5 191 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=107090 $D=1
M21 182 5 192 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=111720 $D=1
M22 193 6 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=107090 $D=1
M23 194 6 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=111720 $D=1
M24 195 193 191 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=107090 $D=1
M25 196 194 192 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=111720 $D=1
M26 189 6 195 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=107090 $D=1
M27 190 6 196 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=111720 $D=1
M28 197 7 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=107090 $D=1
M29 198 7 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=111720 $D=1
M30 199 197 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=107090 $D=1
M31 200 198 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=111720 $D=1
M32 9 7 199 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=107090 $D=1
M33 10 7 200 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=111720 $D=1
M34 201 197 11 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=107090 $D=1
M35 202 198 12 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=111720 $D=1
M36 203 7 201 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=107090 $D=1
M37 204 7 202 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=111720 $D=1
M38 207 197 205 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=107090 $D=1
M39 208 198 206 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=111720 $D=1
M40 195 7 207 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=107090 $D=1
M41 196 7 208 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=111720 $D=1
M42 211 209 207 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=107090 $D=1
M43 212 210 208 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=111720 $D=1
M44 209 13 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=107090 $D=1
M45 210 13 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=111720 $D=1
M46 213 209 201 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=107090 $D=1
M47 214 210 202 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=111720 $D=1
M48 199 13 213 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=107090 $D=1
M49 200 13 214 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=111720 $D=1
M50 215 14 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=107090 $D=1
M51 216 14 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=111720 $D=1
M52 217 215 213 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=107090 $D=1
M53 218 216 214 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=111720 $D=1
M54 211 14 217 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=107090 $D=1
M55 212 14 218 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=111720 $D=1
M56 4 15 219 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=107090 $D=1
M57 8 15 220 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=111720 $D=1
M58 221 16 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=107090 $D=1
M59 222 16 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=111720 $D=1
M60 223 15 217 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=107090 $D=1
M61 224 15 218 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=111720 $D=1
M62 4 223 695 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=107090 $D=1
M63 8 224 696 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=111720 $D=1
M64 225 695 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=107090 $D=1
M65 226 696 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=111720 $D=1
M66 223 219 225 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=107090 $D=1
M67 224 220 226 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=111720 $D=1
M68 225 16 227 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=107090 $D=1
M69 226 16 228 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=111720 $D=1
M70 231 17 225 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=107090 $D=1
M71 232 17 226 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=111720 $D=1
M72 229 17 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=107090 $D=1
M73 230 17 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=111720 $D=1
M74 4 18 233 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=107090 $D=1
M75 8 18 234 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=111720 $D=1
M76 235 19 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=107090 $D=1
M77 236 19 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=111720 $D=1
M78 237 18 217 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=107090 $D=1
M79 238 18 218 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=111720 $D=1
M80 4 237 697 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=107090 $D=1
M81 8 238 698 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=111720 $D=1
M82 239 697 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=107090 $D=1
M83 240 698 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=111720 $D=1
M84 237 233 239 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=107090 $D=1
M85 238 234 240 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=111720 $D=1
M86 239 19 227 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=107090 $D=1
M87 240 19 228 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=111720 $D=1
M88 231 20 239 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=107090 $D=1
M89 232 20 240 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=111720 $D=1
M90 241 20 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=107090 $D=1
M91 242 20 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=111720 $D=1
M92 4 21 243 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=107090 $D=1
M93 8 21 244 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=111720 $D=1
M94 245 22 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=107090 $D=1
M95 246 22 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=111720 $D=1
M96 247 21 217 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=107090 $D=1
M97 248 21 218 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=111720 $D=1
M98 4 247 699 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=107090 $D=1
M99 8 248 700 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=111720 $D=1
M100 249 699 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=107090 $D=1
M101 250 700 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=111720 $D=1
M102 247 243 249 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=107090 $D=1
M103 248 244 250 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=111720 $D=1
M104 249 22 227 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=107090 $D=1
M105 250 22 228 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=111720 $D=1
M106 231 23 249 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=107090 $D=1
M107 232 23 250 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=111720 $D=1
M108 251 23 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=107090 $D=1
M109 252 23 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=111720 $D=1
M110 4 24 253 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=107090 $D=1
M111 8 24 254 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=111720 $D=1
M112 255 25 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=107090 $D=1
M113 256 25 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=111720 $D=1
M114 257 24 217 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=107090 $D=1
M115 258 24 218 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=111720 $D=1
M116 4 257 701 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=107090 $D=1
M117 8 258 702 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=111720 $D=1
M118 259 701 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=107090 $D=1
M119 260 702 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=111720 $D=1
M120 257 253 259 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=107090 $D=1
M121 258 254 260 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=111720 $D=1
M122 259 25 227 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=107090 $D=1
M123 260 25 228 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=111720 $D=1
M124 231 26 259 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=107090 $D=1
M125 232 26 260 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=111720 $D=1
M126 261 26 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=107090 $D=1
M127 262 26 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=111720 $D=1
M128 4 27 263 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=107090 $D=1
M129 8 27 264 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=111720 $D=1
M130 265 28 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=107090 $D=1
M131 266 28 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=111720 $D=1
M132 267 27 217 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=107090 $D=1
M133 268 27 218 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=111720 $D=1
M134 4 267 703 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=107090 $D=1
M135 8 268 704 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=111720 $D=1
M136 269 703 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=107090 $D=1
M137 270 704 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=111720 $D=1
M138 267 263 269 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=107090 $D=1
M139 268 264 270 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=111720 $D=1
M140 269 28 227 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=107090 $D=1
M141 270 28 228 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=111720 $D=1
M142 231 29 269 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=107090 $D=1
M143 232 29 270 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=111720 $D=1
M144 271 29 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=107090 $D=1
M145 272 29 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=111720 $D=1
M146 4 30 273 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=107090 $D=1
M147 8 30 274 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=111720 $D=1
M148 275 31 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=107090 $D=1
M149 276 31 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=111720 $D=1
M150 277 30 217 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=107090 $D=1
M151 278 30 218 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=111720 $D=1
M152 4 277 705 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=107090 $D=1
M153 8 278 706 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=111720 $D=1
M154 279 705 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=107090 $D=1
M155 280 706 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=111720 $D=1
M156 277 273 279 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=107090 $D=1
M157 278 274 280 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=111720 $D=1
M158 279 31 227 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=107090 $D=1
M159 280 31 228 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=111720 $D=1
M160 231 32 279 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=107090 $D=1
M161 232 32 280 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=111720 $D=1
M162 281 32 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=107090 $D=1
M163 282 32 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=111720 $D=1
M164 4 33 283 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=107090 $D=1
M165 8 33 284 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=111720 $D=1
M166 285 34 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=107090 $D=1
M167 286 34 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=111720 $D=1
M168 287 33 217 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=107090 $D=1
M169 288 33 218 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=111720 $D=1
M170 4 287 707 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=107090 $D=1
M171 8 288 708 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=111720 $D=1
M172 289 707 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=107090 $D=1
M173 290 708 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=111720 $D=1
M174 287 283 289 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=107090 $D=1
M175 288 284 290 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=111720 $D=1
M176 289 34 227 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=107090 $D=1
M177 290 34 228 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=111720 $D=1
M178 231 35 289 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=107090 $D=1
M179 232 35 290 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=111720 $D=1
M180 291 35 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=107090 $D=1
M181 292 35 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=111720 $D=1
M182 4 36 293 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=107090 $D=1
M183 8 36 294 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=111720 $D=1
M184 295 37 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=107090 $D=1
M185 296 37 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=111720 $D=1
M186 297 36 217 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=107090 $D=1
M187 298 36 218 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=111720 $D=1
M188 4 297 709 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=107090 $D=1
M189 8 298 710 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=111720 $D=1
M190 299 709 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=107090 $D=1
M191 300 710 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=111720 $D=1
M192 297 293 299 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=107090 $D=1
M193 298 294 300 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=111720 $D=1
M194 299 37 227 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=107090 $D=1
M195 300 37 228 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=111720 $D=1
M196 231 38 299 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=107090 $D=1
M197 232 38 300 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=111720 $D=1
M198 301 38 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=107090 $D=1
M199 302 38 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=111720 $D=1
M200 4 39 303 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=107090 $D=1
M201 8 39 304 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=111720 $D=1
M202 305 40 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=107090 $D=1
M203 306 40 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=111720 $D=1
M204 307 39 217 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=107090 $D=1
M205 308 39 218 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=111720 $D=1
M206 4 307 711 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=107090 $D=1
M207 8 308 712 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=111720 $D=1
M208 309 711 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=107090 $D=1
M209 310 712 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=111720 $D=1
M210 307 303 309 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=107090 $D=1
M211 308 304 310 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=111720 $D=1
M212 309 40 227 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=107090 $D=1
M213 310 40 228 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=111720 $D=1
M214 231 41 309 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=107090 $D=1
M215 232 41 310 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=111720 $D=1
M216 311 41 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=107090 $D=1
M217 312 41 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=111720 $D=1
M218 4 42 313 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=107090 $D=1
M219 8 42 314 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=111720 $D=1
M220 315 43 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=107090 $D=1
M221 316 43 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=111720 $D=1
M222 317 42 217 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=107090 $D=1
M223 318 42 218 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=111720 $D=1
M224 4 317 713 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=107090 $D=1
M225 8 318 714 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=111720 $D=1
M226 319 713 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=107090 $D=1
M227 320 714 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=111720 $D=1
M228 317 313 319 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=107090 $D=1
M229 318 314 320 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=111720 $D=1
M230 319 43 227 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=107090 $D=1
M231 320 43 228 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=111720 $D=1
M232 231 44 319 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=107090 $D=1
M233 232 44 320 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=111720 $D=1
M234 321 44 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=107090 $D=1
M235 322 44 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=111720 $D=1
M236 4 45 323 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=107090 $D=1
M237 8 45 324 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=111720 $D=1
M238 325 46 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=107090 $D=1
M239 326 46 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=111720 $D=1
M240 327 45 217 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=107090 $D=1
M241 328 45 218 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=111720 $D=1
M242 4 327 715 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=107090 $D=1
M243 8 328 716 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=111720 $D=1
M244 329 715 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=107090 $D=1
M245 330 716 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=111720 $D=1
M246 327 323 329 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=107090 $D=1
M247 328 324 330 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=111720 $D=1
M248 329 46 227 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=107090 $D=1
M249 330 46 228 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=111720 $D=1
M250 231 47 329 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=107090 $D=1
M251 232 47 330 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=111720 $D=1
M252 331 47 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=107090 $D=1
M253 332 47 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=111720 $D=1
M254 4 48 333 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=107090 $D=1
M255 8 48 334 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=111720 $D=1
M256 335 49 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=107090 $D=1
M257 336 49 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=111720 $D=1
M258 337 48 217 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=107090 $D=1
M259 338 48 218 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=111720 $D=1
M260 4 337 717 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=107090 $D=1
M261 8 338 718 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=111720 $D=1
M262 339 717 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=107090 $D=1
M263 340 718 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=111720 $D=1
M264 337 333 339 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=107090 $D=1
M265 338 334 340 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=111720 $D=1
M266 339 49 227 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=107090 $D=1
M267 340 49 228 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=111720 $D=1
M268 231 50 339 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=107090 $D=1
M269 232 50 340 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=111720 $D=1
M270 341 50 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=107090 $D=1
M271 342 50 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=111720 $D=1
M272 4 51 343 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=107090 $D=1
M273 8 51 344 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=111720 $D=1
M274 345 52 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=107090 $D=1
M275 346 52 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=111720 $D=1
M276 347 51 217 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=107090 $D=1
M277 348 51 218 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=111720 $D=1
M278 4 347 719 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=107090 $D=1
M279 8 348 720 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=111720 $D=1
M280 349 719 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=107090 $D=1
M281 350 720 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=111720 $D=1
M282 347 343 349 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=107090 $D=1
M283 348 344 350 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=111720 $D=1
M284 349 52 227 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=107090 $D=1
M285 350 52 228 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=111720 $D=1
M286 231 53 349 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=107090 $D=1
M287 232 53 350 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=111720 $D=1
M288 351 53 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=107090 $D=1
M289 352 53 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=111720 $D=1
M290 4 54 353 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=107090 $D=1
M291 8 54 354 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=111720 $D=1
M292 355 55 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=107090 $D=1
M293 356 55 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=111720 $D=1
M294 357 54 217 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=107090 $D=1
M295 358 54 218 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=111720 $D=1
M296 4 357 721 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=107090 $D=1
M297 8 358 722 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=111720 $D=1
M298 359 721 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=107090 $D=1
M299 360 722 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=111720 $D=1
M300 357 353 359 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=107090 $D=1
M301 358 354 360 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=111720 $D=1
M302 359 55 227 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=107090 $D=1
M303 360 55 228 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=111720 $D=1
M304 231 56 359 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=107090 $D=1
M305 232 56 360 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=111720 $D=1
M306 361 56 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=107090 $D=1
M307 362 56 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=111720 $D=1
M308 4 57 363 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=107090 $D=1
M309 8 57 364 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=111720 $D=1
M310 365 58 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=107090 $D=1
M311 366 58 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=111720 $D=1
M312 367 57 217 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=107090 $D=1
M313 368 57 218 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=111720 $D=1
M314 4 367 723 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=107090 $D=1
M315 8 368 724 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=111720 $D=1
M316 369 723 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=107090 $D=1
M317 370 724 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=111720 $D=1
M318 367 363 369 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=107090 $D=1
M319 368 364 370 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=111720 $D=1
M320 369 58 227 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=107090 $D=1
M321 370 58 228 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=111720 $D=1
M322 231 59 369 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=107090 $D=1
M323 232 59 370 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=111720 $D=1
M324 371 59 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=107090 $D=1
M325 372 59 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=111720 $D=1
M326 4 60 373 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=107090 $D=1
M327 8 60 374 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=111720 $D=1
M328 375 61 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=107090 $D=1
M329 376 61 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=111720 $D=1
M330 377 60 217 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=107090 $D=1
M331 378 60 218 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=111720 $D=1
M332 4 377 725 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=107090 $D=1
M333 8 378 726 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=111720 $D=1
M334 379 725 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=107090 $D=1
M335 380 726 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=111720 $D=1
M336 377 373 379 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=107090 $D=1
M337 378 374 380 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=111720 $D=1
M338 379 61 227 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=107090 $D=1
M339 380 61 228 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=111720 $D=1
M340 231 62 379 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=107090 $D=1
M341 232 62 380 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=111720 $D=1
M342 381 62 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=107090 $D=1
M343 382 62 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=111720 $D=1
M344 4 63 383 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=107090 $D=1
M345 8 63 384 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=111720 $D=1
M346 385 64 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=107090 $D=1
M347 386 64 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=111720 $D=1
M348 387 63 217 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=107090 $D=1
M349 388 63 218 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=111720 $D=1
M350 4 387 727 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=107090 $D=1
M351 8 388 728 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=111720 $D=1
M352 389 727 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=107090 $D=1
M353 390 728 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=111720 $D=1
M354 387 383 389 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=107090 $D=1
M355 388 384 390 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=111720 $D=1
M356 389 64 227 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=107090 $D=1
M357 390 64 228 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=111720 $D=1
M358 231 65 389 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=107090 $D=1
M359 232 65 390 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=111720 $D=1
M360 391 65 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=107090 $D=1
M361 392 65 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=111720 $D=1
M362 4 66 393 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=107090 $D=1
M363 8 66 394 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=111720 $D=1
M364 395 67 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=107090 $D=1
M365 396 67 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=111720 $D=1
M366 397 66 217 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=107090 $D=1
M367 398 66 218 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=111720 $D=1
M368 4 397 729 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=107090 $D=1
M369 8 398 730 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=111720 $D=1
M370 399 729 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=107090 $D=1
M371 400 730 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=111720 $D=1
M372 397 393 399 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=107090 $D=1
M373 398 394 400 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=111720 $D=1
M374 399 67 227 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=107090 $D=1
M375 400 67 228 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=111720 $D=1
M376 231 68 399 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=107090 $D=1
M377 232 68 400 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=111720 $D=1
M378 401 68 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=107090 $D=1
M379 402 68 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=111720 $D=1
M380 4 69 403 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=107090 $D=1
M381 8 69 404 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=111720 $D=1
M382 405 70 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=107090 $D=1
M383 406 70 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=111720 $D=1
M384 407 69 217 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=107090 $D=1
M385 408 69 218 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=111720 $D=1
M386 4 407 731 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=107090 $D=1
M387 8 408 732 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=111720 $D=1
M388 409 731 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=107090 $D=1
M389 410 732 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=111720 $D=1
M390 407 403 409 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=107090 $D=1
M391 408 404 410 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=111720 $D=1
M392 409 70 227 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=107090 $D=1
M393 410 70 228 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=111720 $D=1
M394 231 71 409 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=107090 $D=1
M395 232 71 410 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=111720 $D=1
M396 411 71 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=107090 $D=1
M397 412 71 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=111720 $D=1
M398 4 72 413 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=107090 $D=1
M399 8 72 414 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=111720 $D=1
M400 415 73 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=107090 $D=1
M401 416 73 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=111720 $D=1
M402 417 72 217 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=107090 $D=1
M403 418 72 218 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=111720 $D=1
M404 4 417 733 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=107090 $D=1
M405 8 418 734 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=111720 $D=1
M406 419 733 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=107090 $D=1
M407 420 734 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=111720 $D=1
M408 417 413 419 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=107090 $D=1
M409 418 414 420 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=111720 $D=1
M410 419 73 227 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=107090 $D=1
M411 420 73 228 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=111720 $D=1
M412 231 74 419 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=107090 $D=1
M413 232 74 420 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=111720 $D=1
M414 421 74 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=107090 $D=1
M415 422 74 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=111720 $D=1
M416 4 75 423 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=107090 $D=1
M417 8 75 424 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=111720 $D=1
M418 425 76 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=107090 $D=1
M419 426 76 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=111720 $D=1
M420 427 75 217 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=107090 $D=1
M421 428 75 218 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=111720 $D=1
M422 4 427 735 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=107090 $D=1
M423 8 428 736 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=111720 $D=1
M424 429 735 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=107090 $D=1
M425 430 736 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=111720 $D=1
M426 427 423 429 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=107090 $D=1
M427 428 424 430 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=111720 $D=1
M428 429 76 227 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=107090 $D=1
M429 430 76 228 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=111720 $D=1
M430 231 77 429 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=107090 $D=1
M431 232 77 430 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=111720 $D=1
M432 431 77 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=107090 $D=1
M433 432 77 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=111720 $D=1
M434 4 78 433 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=107090 $D=1
M435 8 78 434 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=111720 $D=1
M436 435 79 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=107090 $D=1
M437 436 79 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=111720 $D=1
M438 437 78 217 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=107090 $D=1
M439 438 78 218 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=111720 $D=1
M440 4 437 737 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=107090 $D=1
M441 8 438 738 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=111720 $D=1
M442 439 737 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=107090 $D=1
M443 440 738 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=111720 $D=1
M444 437 433 439 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=107090 $D=1
M445 438 434 440 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=111720 $D=1
M446 439 79 227 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=107090 $D=1
M447 440 79 228 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=111720 $D=1
M448 231 80 439 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=107090 $D=1
M449 232 80 440 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=111720 $D=1
M450 441 80 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=107090 $D=1
M451 442 80 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=111720 $D=1
M452 4 81 443 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=107090 $D=1
M453 8 81 444 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=111720 $D=1
M454 445 82 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=107090 $D=1
M455 446 82 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=111720 $D=1
M456 447 81 217 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=107090 $D=1
M457 448 81 218 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=111720 $D=1
M458 4 447 739 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=107090 $D=1
M459 8 448 740 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=111720 $D=1
M460 449 739 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=107090 $D=1
M461 450 740 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=111720 $D=1
M462 447 443 449 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=107090 $D=1
M463 448 444 450 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=111720 $D=1
M464 449 82 227 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=107090 $D=1
M465 450 82 228 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=111720 $D=1
M466 231 83 449 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=107090 $D=1
M467 232 83 450 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=111720 $D=1
M468 451 83 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=107090 $D=1
M469 452 83 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=111720 $D=1
M470 4 84 453 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=107090 $D=1
M471 8 84 454 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=111720 $D=1
M472 455 85 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=107090 $D=1
M473 456 85 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=111720 $D=1
M474 457 84 217 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=107090 $D=1
M475 458 84 218 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=111720 $D=1
M476 4 457 741 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=107090 $D=1
M477 8 458 742 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=111720 $D=1
M478 459 741 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=107090 $D=1
M479 460 742 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=111720 $D=1
M480 457 453 459 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=107090 $D=1
M481 458 454 460 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=111720 $D=1
M482 459 85 227 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=107090 $D=1
M483 460 85 228 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=111720 $D=1
M484 231 86 459 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=107090 $D=1
M485 232 86 460 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=111720 $D=1
M486 461 86 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=107090 $D=1
M487 462 86 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=111720 $D=1
M488 4 87 463 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=107090 $D=1
M489 8 87 464 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=111720 $D=1
M490 465 88 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=107090 $D=1
M491 466 88 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=111720 $D=1
M492 467 87 217 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=107090 $D=1
M493 468 87 218 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=111720 $D=1
M494 4 467 743 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=107090 $D=1
M495 8 468 744 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=111720 $D=1
M496 469 743 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=107090 $D=1
M497 470 744 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=111720 $D=1
M498 467 463 469 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=107090 $D=1
M499 468 464 470 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=111720 $D=1
M500 469 88 227 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=107090 $D=1
M501 470 88 228 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=111720 $D=1
M502 231 89 469 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=107090 $D=1
M503 232 89 470 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=111720 $D=1
M504 471 89 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=107090 $D=1
M505 472 89 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=111720 $D=1
M506 4 90 473 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=107090 $D=1
M507 8 90 474 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=111720 $D=1
M508 475 91 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=107090 $D=1
M509 476 91 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=111720 $D=1
M510 477 90 217 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=107090 $D=1
M511 478 90 218 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=111720 $D=1
M512 4 477 745 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=107090 $D=1
M513 8 478 746 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=111720 $D=1
M514 479 745 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=107090 $D=1
M515 480 746 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=111720 $D=1
M516 477 473 479 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=107090 $D=1
M517 478 474 480 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=111720 $D=1
M518 479 91 227 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=107090 $D=1
M519 480 91 228 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=111720 $D=1
M520 231 92 479 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=107090 $D=1
M521 232 92 480 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=111720 $D=1
M522 481 92 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=107090 $D=1
M523 482 92 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=111720 $D=1
M524 4 93 483 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=107090 $D=1
M525 8 93 484 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=111720 $D=1
M526 485 94 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=107090 $D=1
M527 486 94 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=111720 $D=1
M528 487 93 217 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=107090 $D=1
M529 488 93 218 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=111720 $D=1
M530 4 487 747 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=107090 $D=1
M531 8 488 748 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=111720 $D=1
M532 489 747 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=107090 $D=1
M533 490 748 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=111720 $D=1
M534 487 483 489 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=107090 $D=1
M535 488 484 490 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=111720 $D=1
M536 489 94 227 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=107090 $D=1
M537 490 94 228 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=111720 $D=1
M538 231 95 489 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=107090 $D=1
M539 232 95 490 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=111720 $D=1
M540 491 95 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=107090 $D=1
M541 492 95 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=111720 $D=1
M542 4 96 493 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=107090 $D=1
M543 8 96 494 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=111720 $D=1
M544 495 97 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=107090 $D=1
M545 496 97 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=111720 $D=1
M546 497 96 217 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=107090 $D=1
M547 498 96 218 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=111720 $D=1
M548 4 497 749 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=107090 $D=1
M549 8 498 750 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=111720 $D=1
M550 499 749 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=107090 $D=1
M551 500 750 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=111720 $D=1
M552 497 493 499 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=107090 $D=1
M553 498 494 500 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=111720 $D=1
M554 499 97 227 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=107090 $D=1
M555 500 97 228 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=111720 $D=1
M556 231 98 499 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=107090 $D=1
M557 232 98 500 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=111720 $D=1
M558 501 98 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=107090 $D=1
M559 502 98 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=111720 $D=1
M560 4 99 503 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=107090 $D=1
M561 8 99 504 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=111720 $D=1
M562 505 100 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=107090 $D=1
M563 506 100 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=111720 $D=1
M564 507 99 217 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=107090 $D=1
M565 508 99 218 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=111720 $D=1
M566 4 507 751 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=107090 $D=1
M567 8 508 752 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=111720 $D=1
M568 509 751 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=107090 $D=1
M569 510 752 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=111720 $D=1
M570 507 503 509 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=107090 $D=1
M571 508 504 510 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=111720 $D=1
M572 509 100 227 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=107090 $D=1
M573 510 100 228 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=111720 $D=1
M574 231 101 509 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=107090 $D=1
M575 232 101 510 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=111720 $D=1
M576 511 101 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=107090 $D=1
M577 512 101 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=111720 $D=1
M578 4 102 513 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=107090 $D=1
M579 8 102 514 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=111720 $D=1
M580 515 103 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=107090 $D=1
M581 516 103 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=111720 $D=1
M582 517 102 217 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=107090 $D=1
M583 518 102 218 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=111720 $D=1
M584 4 517 753 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=107090 $D=1
M585 8 518 754 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=111720 $D=1
M586 519 753 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=107090 $D=1
M587 520 754 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=111720 $D=1
M588 517 513 519 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=107090 $D=1
M589 518 514 520 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=111720 $D=1
M590 519 103 227 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=107090 $D=1
M591 520 103 228 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=111720 $D=1
M592 231 104 519 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=107090 $D=1
M593 232 104 520 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=111720 $D=1
M594 521 104 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=107090 $D=1
M595 522 104 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=111720 $D=1
M596 4 105 523 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=107090 $D=1
M597 8 105 524 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=111720 $D=1
M598 525 106 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=107090 $D=1
M599 526 106 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=111720 $D=1
M600 527 105 217 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=107090 $D=1
M601 528 105 218 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=111720 $D=1
M602 4 527 755 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=107090 $D=1
M603 8 528 756 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=111720 $D=1
M604 529 755 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=107090 $D=1
M605 530 756 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=111720 $D=1
M606 527 523 529 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=107090 $D=1
M607 528 524 530 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=111720 $D=1
M608 529 106 227 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=107090 $D=1
M609 530 106 228 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=111720 $D=1
M610 231 107 529 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=107090 $D=1
M611 232 107 530 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=111720 $D=1
M612 531 107 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=107090 $D=1
M613 532 107 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=111720 $D=1
M614 4 108 533 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=107090 $D=1
M615 8 108 534 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=111720 $D=1
M616 535 109 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=107090 $D=1
M617 536 109 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=111720 $D=1
M618 4 109 227 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=107090 $D=1
M619 8 109 228 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=111720 $D=1
M620 231 108 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=107090 $D=1
M621 232 108 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=111720 $D=1
M622 4 539 537 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=107090 $D=1
M623 8 540 538 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=111720 $D=1
M624 539 110 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=107090 $D=1
M625 540 110 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=111720 $D=1
M626 757 227 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=107090 $D=1
M627 758 228 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=111720 $D=1
M628 541 537 757 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=107090 $D=1
M629 542 538 758 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=111720 $D=1
M630 4 541 543 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=107090 $D=1
M631 8 542 544 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=111720 $D=1
M632 759 543 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=107090 $D=1
M633 760 544 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=111720 $D=1
M634 541 539 759 4 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=107090 $D=1
M635 542 540 760 8 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=111720 $D=1
M636 4 547 545 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=107090 $D=1
M637 8 548 546 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=111720 $D=1
M638 547 110 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=107090 $D=1
M639 548 110 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=111720 $D=1
M640 761 231 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=107090 $D=1
M641 762 232 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=111720 $D=1
M642 549 545 761 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=107090 $D=1
M643 550 546 762 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=111720 $D=1
M644 4 549 111 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=107090 $D=1
M645 8 550 112 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=111720 $D=1
M646 763 111 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=107090 $D=1
M647 764 112 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=111720 $D=1
M648 549 547 763 4 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=107090 $D=1
M649 550 548 764 8 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=111720 $D=1
M650 551 113 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=107090 $D=1
M651 552 113 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=111720 $D=1
M652 553 551 543 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=107090 $D=1
M653 554 552 544 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=111720 $D=1
M654 114 113 553 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=107090 $D=1
M655 115 113 554 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=111720 $D=1
M656 555 116 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=107090 $D=1
M657 556 116 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=111720 $D=1
M658 557 555 111 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=107090 $D=1
M659 558 556 112 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=111720 $D=1
M660 765 116 557 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=107090 $D=1
M661 766 116 558 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=111720 $D=1
M662 4 111 765 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=107090 $D=1
M663 8 112 766 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=111720 $D=1
M664 559 117 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=107090 $D=1
M665 560 117 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=111720 $D=1
M666 561 559 557 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=107090 $D=1
M667 562 560 558 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=111720 $D=1
M668 9 117 561 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=107090 $D=1
M669 10 117 562 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=111720 $D=1
M670 564 563 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=107090 $D=1
M671 565 118 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=111720 $D=1
M672 4 568 566 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=107090 $D=1
M673 8 569 567 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=111720 $D=1
M674 570 553 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=107090 $D=1
M675 571 554 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=111720 $D=1
M676 568 570 563 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=107090 $D=1
M677 569 571 118 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=111720 $D=1
M678 564 553 568 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=107090 $D=1
M679 565 554 569 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=111720 $D=1
M680 572 566 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=107090 $D=1
M681 573 567 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=111720 $D=1
M682 574 572 561 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=107090 $D=1
M683 563 573 562 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=111720 $D=1
M684 553 566 574 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=107090 $D=1
M685 554 567 563 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=111720 $D=1
M686 575 574 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=107090 $D=1
M687 576 563 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=111720 $D=1
M688 577 566 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=107090 $D=1
M689 578 567 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=111720 $D=1
M690 579 577 575 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=107090 $D=1
M691 580 578 576 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=111720 $D=1
M692 561 566 579 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=107090 $D=1
M693 562 567 580 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=111720 $D=1
M694 581 553 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=107090 $D=1
M695 582 554 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=111720 $D=1
M696 4 561 581 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=107090 $D=1
M697 8 562 582 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=111720 $D=1
M698 583 579 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=107090 $D=1
M699 584 580 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=111720 $D=1
M700 796 553 4 4 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=107090 $D=1
M701 797 554 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=111720 $D=1
M702 585 561 796 4 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=107090 $D=1
M703 586 562 797 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=111720 $D=1
M704 798 553 4 4 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=107090 $D=1
M705 799 554 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=111720 $D=1
M706 587 561 798 4 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=107090 $D=1
M707 588 562 799 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=111720 $D=1
M708 591 553 589 4 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=107090 $D=1
M709 592 554 590 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=111720 $D=1
M710 589 561 591 4 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=107090 $D=1
M711 590 562 592 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=111720 $D=1
M712 4 587 589 4 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=107090 $D=1
M713 8 588 590 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=111720 $D=1
M714 593 119 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=107090 $D=1
M715 594 119 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=111720 $D=1
M716 595 593 581 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=107090 $D=1
M717 596 594 582 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=111720 $D=1
M718 585 119 595 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=107090 $D=1
M719 586 119 596 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=111720 $D=1
M720 597 593 583 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=107090 $D=1
M721 598 594 584 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=111720 $D=1
M722 591 119 597 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=107090 $D=1
M723 592 119 598 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=111720 $D=1
M724 599 120 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=107090 $D=1
M725 600 120 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=111720 $D=1
M726 601 599 597 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=107090 $D=1
M727 602 600 598 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=111720 $D=1
M728 595 120 601 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=107090 $D=1
M729 596 120 602 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=111720 $D=1
M730 11 601 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=107090 $D=1
M731 12 602 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=111720 $D=1
M732 603 121 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=107090 $D=1
M733 604 121 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=111720 $D=1
M734 605 603 122 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=107090 $D=1
M735 606 604 123 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=111720 $D=1
M736 124 121 605 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=107090 $D=1
M737 125 121 606 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=111720 $D=1
M738 607 121 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=107090 $D=1
M739 608 121 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=111720 $D=1
M740 613 607 127 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=107090 $D=1
M741 614 608 129 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=111720 $D=1
M742 130 121 613 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=107090 $D=1
M743 128 121 614 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=111720 $D=1
M744 615 121 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=107090 $D=1
M745 616 121 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=111720 $D=1
M746 133 615 131 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=107090 $D=1
M747 133 616 132 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=111720 $D=1
M748 134 121 133 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=107090 $D=1
M749 135 121 133 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=111720 $D=1
M750 617 121 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=107090 $D=1
M751 618 121 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=111720 $D=1
M752 619 617 136 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=107090 $D=1
M753 620 618 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=111720 $D=1
M754 137 121 619 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=107090 $D=1
M755 138 121 620 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=111720 $D=1
M756 621 121 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=107090 $D=1
M757 622 121 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=111720 $D=1
M758 623 621 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=107090 $D=1
M759 624 622 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=111720 $D=1
M760 139 121 623 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=107090 $D=1
M761 140 121 624 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=111720 $D=1
M762 4 553 778 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=107090 $D=1
M763 8 554 779 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=111720 $D=1
M764 125 778 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=107090 $D=1
M765 122 779 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=111720 $D=1
M766 625 141 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=107090 $D=1
M767 626 141 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=111720 $D=1
M768 143 625 125 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=107090 $D=1
M769 144 626 122 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=111720 $D=1
M770 605 141 143 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=107090 $D=1
M771 606 141 144 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=111720 $D=1
M772 627 145 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=107090 $D=1
M773 628 145 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=111720 $D=1
M774 126 627 143 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=107090 $D=1
M775 146 628 144 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=111720 $D=1
M776 613 145 126 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=107090 $D=1
M777 614 145 146 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=111720 $D=1
M778 629 147 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=107090 $D=1
M779 630 147 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=111720 $D=1
M780 142 629 126 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=107090 $D=1
M781 148 630 146 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=111720 $D=1
M782 133 147 142 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=107090 $D=1
M783 133 147 148 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=111720 $D=1
M784 631 149 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=107090 $D=1
M785 632 149 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=111720 $D=1
M786 150 631 142 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=107090 $D=1
M787 151 632 148 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=111720 $D=1
M788 619 149 150 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=107090 $D=1
M789 620 149 151 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=111720 $D=1
M790 633 152 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=107090 $D=1
M791 634 152 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=111720 $D=1
M792 203 633 150 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=107090 $D=1
M793 204 634 151 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=111720 $D=1
M794 623 152 203 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=107090 $D=1
M795 624 152 204 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=111720 $D=1
M796 635 153 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=107090 $D=1
M797 636 153 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=111720 $D=1
M798 637 635 111 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=107090 $D=1
M799 638 636 112 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=111720 $D=1
M800 9 153 637 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=107090 $D=1
M801 10 153 638 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=111720 $D=1
M802 800 543 4 4 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=107090 $D=1
M803 801 544 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=111720 $D=1
M804 639 637 800 4 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=107090 $D=1
M805 640 638 801 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=111720 $D=1
M806 643 543 641 4 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=107090 $D=1
M807 644 544 642 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=111720 $D=1
M808 641 637 643 4 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=107090 $D=1
M809 642 638 644 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=111720 $D=1
M810 4 639 641 4 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=107090 $D=1
M811 8 640 642 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=111720 $D=1
M812 802 645 4 4 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=107090 $D=1
M813 803 646 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=111720 $D=1
M814 780 643 802 4 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=107090 $D=1
M815 781 644 803 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=111720 $D=1
M816 646 780 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=107090 $D=1
M817 154 781 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=111720 $D=1
M818 647 543 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=107090 $D=1
M819 648 544 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=111720 $D=1
M820 4 649 647 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=107090 $D=1
M821 8 650 648 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=111720 $D=1
M822 649 637 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=107090 $D=1
M823 650 638 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=111720 $D=1
M824 804 647 4 4 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=107090 $D=1
M825 805 648 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=111720 $D=1
M826 651 645 804 4 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=107090 $D=1
M827 652 646 805 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=111720 $D=1
M828 654 155 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=107090 $D=1
M829 655 653 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=111720 $D=1
M830 806 651 4 4 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=107090 $D=1
M831 807 652 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=111720 $D=1
M832 653 654 806 4 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=107090 $D=1
M833 156 655 807 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=111720 $D=1
M834 657 656 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=107090 $D=1
M835 658 157 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=111720 $D=1
M836 4 661 659 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=107090 $D=1
M837 8 662 660 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=111720 $D=1
M838 663 114 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=107090 $D=1
M839 664 115 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=111720 $D=1
M840 661 663 656 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=107090 $D=1
M841 662 664 157 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=111720 $D=1
M842 657 114 661 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=107090 $D=1
M843 658 115 662 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=111720 $D=1
M844 665 659 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=107090 $D=1
M845 666 660 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=111720 $D=1
M846 158 665 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=107090 $D=1
M847 656 666 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=111720 $D=1
M848 114 659 158 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=107090 $D=1
M849 115 660 656 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=111720 $D=1
M850 667 158 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=107090 $D=1
M851 668 656 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=111720 $D=1
M852 669 659 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=107090 $D=1
M853 670 660 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=111720 $D=1
M854 205 669 667 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=107090 $D=1
M855 206 670 668 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=111720 $D=1
M856 4 659 205 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=107090 $D=1
M857 8 660 206 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=111720 $D=1
M858 671 159 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=107090 $D=1
M859 672 159 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=111720 $D=1
M860 673 671 205 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=107090 $D=1
M861 674 672 206 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=111720 $D=1
M862 11 159 673 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=107090 $D=1
M863 12 159 674 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=111720 $D=1
M864 675 160 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=107090 $D=1
M865 676 160 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=111720 $D=1
M866 160 675 673 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=107090 $D=1
M867 160 676 674 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=111720 $D=1
M868 4 160 160 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=107090 $D=1
M869 8 160 160 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=111720 $D=1
M870 677 110 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=107090 $D=1
M871 678 110 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=111720 $D=1
M872 4 677 679 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=107090 $D=1
M873 8 678 680 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=111720 $D=1
M874 681 110 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=107090 $D=1
M875 682 110 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=111720 $D=1
M876 683 677 160 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=107090 $D=1
M877 684 678 160 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=111720 $D=1
M878 4 683 782 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=107090 $D=1
M879 8 684 783 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=111720 $D=1
M880 685 782 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=107090 $D=1
M881 686 783 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=111720 $D=1
M882 683 679 685 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=107090 $D=1
M883 684 680 686 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=111720 $D=1
M884 687 110 685 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=107090 $D=1
M885 688 110 686 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=111720 $D=1
M886 4 691 689 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=107090 $D=1
M887 8 692 690 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=111720 $D=1
M888 691 110 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=107090 $D=1
M889 692 110 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=111720 $D=1
M890 784 687 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=107090 $D=1
M891 785 688 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=111720 $D=1
M892 693 689 784 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=107090 $D=1
M893 694 690 785 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=111720 $D=1
M894 4 693 114 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=107090 $D=1
M895 8 694 115 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=111720 $D=1
M896 786 114 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=107090 $D=1
M897 787 115 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=111720 $D=1
M898 693 691 786 4 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=107090 $D=1
M899 694 692 787 8 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=111720 $D=1
M900 179 1 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=108340 $D=0
M901 180 1 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=112970 $D=0
M902 181 1 2 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=108340 $D=0
M903 182 1 3 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=112970 $D=0
M904 4 179 181 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=108340 $D=0
M905 8 180 182 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=112970 $D=0
M906 183 1 3 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=108340 $D=0
M907 184 1 3 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=112970 $D=0
M908 2 179 183 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=108340 $D=0
M909 3 180 184 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=112970 $D=0
M910 185 1 4 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=108340 $D=0
M911 186 1 3 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=112970 $D=0
M912 2 179 185 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=108340 $D=0
M913 3 180 186 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=112970 $D=0
M914 189 5 185 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=108340 $D=0
M915 190 5 186 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=112970 $D=0
M916 187 5 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=108340 $D=0
M917 188 5 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=112970 $D=0
M918 191 5 183 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=108340 $D=0
M919 192 5 184 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=112970 $D=0
M920 181 187 191 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=108340 $D=0
M921 182 188 192 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=112970 $D=0
M922 193 6 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=108340 $D=0
M923 194 6 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=112970 $D=0
M924 195 6 191 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=108340 $D=0
M925 196 6 192 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=112970 $D=0
M926 189 193 195 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=108340 $D=0
M927 190 194 196 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=112970 $D=0
M928 197 7 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=108340 $D=0
M929 198 7 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=112970 $D=0
M930 199 7 4 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=108340 $D=0
M931 200 7 8 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=112970 $D=0
M932 9 197 199 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=108340 $D=0
M933 10 198 200 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=112970 $D=0
M934 201 7 11 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=108340 $D=0
M935 202 7 12 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=112970 $D=0
M936 203 197 201 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=108340 $D=0
M937 204 198 202 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=112970 $D=0
M938 207 7 205 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=108340 $D=0
M939 208 7 206 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=112970 $D=0
M940 195 197 207 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=108340 $D=0
M941 196 198 208 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=112970 $D=0
M942 211 13 207 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=108340 $D=0
M943 212 13 208 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=112970 $D=0
M944 209 13 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=108340 $D=0
M945 210 13 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=112970 $D=0
M946 213 13 201 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=108340 $D=0
M947 214 13 202 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=112970 $D=0
M948 199 209 213 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=108340 $D=0
M949 200 210 214 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=112970 $D=0
M950 215 14 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=108340 $D=0
M951 216 14 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=112970 $D=0
M952 217 14 213 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=108340 $D=0
M953 218 14 214 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=112970 $D=0
M954 211 215 217 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=108340 $D=0
M955 212 216 218 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=112970 $D=0
M956 161 15 219 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=108340 $D=0
M957 162 15 220 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=112970 $D=0
M958 221 16 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=108340 $D=0
M959 222 16 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=112970 $D=0
M960 223 219 217 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=108340 $D=0
M961 224 220 218 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=112970 $D=0
M962 161 223 695 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=108340 $D=0
M963 162 224 696 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=112970 $D=0
M964 225 695 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=108340 $D=0
M965 226 696 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=112970 $D=0
M966 223 15 225 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=108340 $D=0
M967 224 15 226 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=112970 $D=0
M968 225 221 227 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=108340 $D=0
M969 226 222 228 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=112970 $D=0
M970 231 229 225 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=108340 $D=0
M971 232 230 226 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=112970 $D=0
M972 229 17 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=108340 $D=0
M973 230 17 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=112970 $D=0
M974 161 18 233 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=108340 $D=0
M975 162 18 234 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=112970 $D=0
M976 235 19 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=108340 $D=0
M977 236 19 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=112970 $D=0
M978 237 233 217 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=108340 $D=0
M979 238 234 218 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=112970 $D=0
M980 161 237 697 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=108340 $D=0
M981 162 238 698 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=112970 $D=0
M982 239 697 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=108340 $D=0
M983 240 698 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=112970 $D=0
M984 237 18 239 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=108340 $D=0
M985 238 18 240 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=112970 $D=0
M986 239 235 227 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=108340 $D=0
M987 240 236 228 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=112970 $D=0
M988 231 241 239 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=108340 $D=0
M989 232 242 240 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=112970 $D=0
M990 241 20 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=108340 $D=0
M991 242 20 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=112970 $D=0
M992 161 21 243 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=108340 $D=0
M993 162 21 244 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=112970 $D=0
M994 245 22 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=108340 $D=0
M995 246 22 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=112970 $D=0
M996 247 243 217 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=108340 $D=0
M997 248 244 218 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=112970 $D=0
M998 161 247 699 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=108340 $D=0
M999 162 248 700 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=112970 $D=0
M1000 249 699 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=108340 $D=0
M1001 250 700 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=112970 $D=0
M1002 247 21 249 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=108340 $D=0
M1003 248 21 250 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=112970 $D=0
M1004 249 245 227 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=108340 $D=0
M1005 250 246 228 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=112970 $D=0
M1006 231 251 249 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=108340 $D=0
M1007 232 252 250 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=112970 $D=0
M1008 251 23 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=108340 $D=0
M1009 252 23 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=112970 $D=0
M1010 161 24 253 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=108340 $D=0
M1011 162 24 254 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=112970 $D=0
M1012 255 25 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=108340 $D=0
M1013 256 25 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=112970 $D=0
M1014 257 253 217 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=108340 $D=0
M1015 258 254 218 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=112970 $D=0
M1016 161 257 701 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=108340 $D=0
M1017 162 258 702 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=112970 $D=0
M1018 259 701 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=108340 $D=0
M1019 260 702 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=112970 $D=0
M1020 257 24 259 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=108340 $D=0
M1021 258 24 260 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=112970 $D=0
M1022 259 255 227 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=108340 $D=0
M1023 260 256 228 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=112970 $D=0
M1024 231 261 259 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=108340 $D=0
M1025 232 262 260 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=112970 $D=0
M1026 261 26 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=108340 $D=0
M1027 262 26 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=112970 $D=0
M1028 161 27 263 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=108340 $D=0
M1029 162 27 264 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=112970 $D=0
M1030 265 28 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=108340 $D=0
M1031 266 28 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=112970 $D=0
M1032 267 263 217 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=108340 $D=0
M1033 268 264 218 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=112970 $D=0
M1034 161 267 703 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=108340 $D=0
M1035 162 268 704 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=112970 $D=0
M1036 269 703 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=108340 $D=0
M1037 270 704 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=112970 $D=0
M1038 267 27 269 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=108340 $D=0
M1039 268 27 270 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=112970 $D=0
M1040 269 265 227 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=108340 $D=0
M1041 270 266 228 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=112970 $D=0
M1042 231 271 269 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=108340 $D=0
M1043 232 272 270 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=112970 $D=0
M1044 271 29 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=108340 $D=0
M1045 272 29 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=112970 $D=0
M1046 161 30 273 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=108340 $D=0
M1047 162 30 274 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=112970 $D=0
M1048 275 31 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=108340 $D=0
M1049 276 31 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=112970 $D=0
M1050 277 273 217 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=108340 $D=0
M1051 278 274 218 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=112970 $D=0
M1052 161 277 705 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=108340 $D=0
M1053 162 278 706 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=112970 $D=0
M1054 279 705 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=108340 $D=0
M1055 280 706 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=112970 $D=0
M1056 277 30 279 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=108340 $D=0
M1057 278 30 280 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=112970 $D=0
M1058 279 275 227 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=108340 $D=0
M1059 280 276 228 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=112970 $D=0
M1060 231 281 279 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=108340 $D=0
M1061 232 282 280 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=112970 $D=0
M1062 281 32 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=108340 $D=0
M1063 282 32 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=112970 $D=0
M1064 161 33 283 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=108340 $D=0
M1065 162 33 284 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=112970 $D=0
M1066 285 34 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=108340 $D=0
M1067 286 34 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=112970 $D=0
M1068 287 283 217 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=108340 $D=0
M1069 288 284 218 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=112970 $D=0
M1070 161 287 707 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=108340 $D=0
M1071 162 288 708 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=112970 $D=0
M1072 289 707 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=108340 $D=0
M1073 290 708 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=112970 $D=0
M1074 287 33 289 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=108340 $D=0
M1075 288 33 290 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=112970 $D=0
M1076 289 285 227 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=108340 $D=0
M1077 290 286 228 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=112970 $D=0
M1078 231 291 289 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=108340 $D=0
M1079 232 292 290 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=112970 $D=0
M1080 291 35 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=108340 $D=0
M1081 292 35 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=112970 $D=0
M1082 161 36 293 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=108340 $D=0
M1083 162 36 294 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=112970 $D=0
M1084 295 37 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=108340 $D=0
M1085 296 37 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=112970 $D=0
M1086 297 293 217 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=108340 $D=0
M1087 298 294 218 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=112970 $D=0
M1088 161 297 709 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=108340 $D=0
M1089 162 298 710 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=112970 $D=0
M1090 299 709 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=108340 $D=0
M1091 300 710 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=112970 $D=0
M1092 297 36 299 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=108340 $D=0
M1093 298 36 300 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=112970 $D=0
M1094 299 295 227 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=108340 $D=0
M1095 300 296 228 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=112970 $D=0
M1096 231 301 299 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=108340 $D=0
M1097 232 302 300 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=112970 $D=0
M1098 301 38 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=108340 $D=0
M1099 302 38 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=112970 $D=0
M1100 161 39 303 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=108340 $D=0
M1101 162 39 304 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=112970 $D=0
M1102 305 40 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=108340 $D=0
M1103 306 40 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=112970 $D=0
M1104 307 303 217 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=108340 $D=0
M1105 308 304 218 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=112970 $D=0
M1106 161 307 711 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=108340 $D=0
M1107 162 308 712 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=112970 $D=0
M1108 309 711 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=108340 $D=0
M1109 310 712 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=112970 $D=0
M1110 307 39 309 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=108340 $D=0
M1111 308 39 310 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=112970 $D=0
M1112 309 305 227 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=108340 $D=0
M1113 310 306 228 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=112970 $D=0
M1114 231 311 309 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=108340 $D=0
M1115 232 312 310 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=112970 $D=0
M1116 311 41 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=108340 $D=0
M1117 312 41 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=112970 $D=0
M1118 161 42 313 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=108340 $D=0
M1119 162 42 314 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=112970 $D=0
M1120 315 43 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=108340 $D=0
M1121 316 43 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=112970 $D=0
M1122 317 313 217 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=108340 $D=0
M1123 318 314 218 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=112970 $D=0
M1124 161 317 713 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=108340 $D=0
M1125 162 318 714 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=112970 $D=0
M1126 319 713 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=108340 $D=0
M1127 320 714 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=112970 $D=0
M1128 317 42 319 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=108340 $D=0
M1129 318 42 320 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=112970 $D=0
M1130 319 315 227 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=108340 $D=0
M1131 320 316 228 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=112970 $D=0
M1132 231 321 319 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=108340 $D=0
M1133 232 322 320 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=112970 $D=0
M1134 321 44 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=108340 $D=0
M1135 322 44 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=112970 $D=0
M1136 161 45 323 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=108340 $D=0
M1137 162 45 324 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=112970 $D=0
M1138 325 46 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=108340 $D=0
M1139 326 46 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=112970 $D=0
M1140 327 323 217 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=108340 $D=0
M1141 328 324 218 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=112970 $D=0
M1142 161 327 715 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=108340 $D=0
M1143 162 328 716 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=112970 $D=0
M1144 329 715 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=108340 $D=0
M1145 330 716 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=112970 $D=0
M1146 327 45 329 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=108340 $D=0
M1147 328 45 330 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=112970 $D=0
M1148 329 325 227 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=108340 $D=0
M1149 330 326 228 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=112970 $D=0
M1150 231 331 329 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=108340 $D=0
M1151 232 332 330 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=112970 $D=0
M1152 331 47 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=108340 $D=0
M1153 332 47 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=112970 $D=0
M1154 161 48 333 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=108340 $D=0
M1155 162 48 334 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=112970 $D=0
M1156 335 49 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=108340 $D=0
M1157 336 49 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=112970 $D=0
M1158 337 333 217 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=108340 $D=0
M1159 338 334 218 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=112970 $D=0
M1160 161 337 717 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=108340 $D=0
M1161 162 338 718 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=112970 $D=0
M1162 339 717 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=108340 $D=0
M1163 340 718 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=112970 $D=0
M1164 337 48 339 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=108340 $D=0
M1165 338 48 340 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=112970 $D=0
M1166 339 335 227 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=108340 $D=0
M1167 340 336 228 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=112970 $D=0
M1168 231 341 339 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=108340 $D=0
M1169 232 342 340 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=112970 $D=0
M1170 341 50 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=108340 $D=0
M1171 342 50 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=112970 $D=0
M1172 161 51 343 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=108340 $D=0
M1173 162 51 344 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=112970 $D=0
M1174 345 52 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=108340 $D=0
M1175 346 52 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=112970 $D=0
M1176 347 343 217 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=108340 $D=0
M1177 348 344 218 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=112970 $D=0
M1178 161 347 719 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=108340 $D=0
M1179 162 348 720 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=112970 $D=0
M1180 349 719 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=108340 $D=0
M1181 350 720 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=112970 $D=0
M1182 347 51 349 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=108340 $D=0
M1183 348 51 350 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=112970 $D=0
M1184 349 345 227 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=108340 $D=0
M1185 350 346 228 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=112970 $D=0
M1186 231 351 349 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=108340 $D=0
M1187 232 352 350 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=112970 $D=0
M1188 351 53 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=108340 $D=0
M1189 352 53 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=112970 $D=0
M1190 161 54 353 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=108340 $D=0
M1191 162 54 354 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=112970 $D=0
M1192 355 55 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=108340 $D=0
M1193 356 55 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=112970 $D=0
M1194 357 353 217 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=108340 $D=0
M1195 358 354 218 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=112970 $D=0
M1196 161 357 721 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=108340 $D=0
M1197 162 358 722 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=112970 $D=0
M1198 359 721 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=108340 $D=0
M1199 360 722 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=112970 $D=0
M1200 357 54 359 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=108340 $D=0
M1201 358 54 360 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=112970 $D=0
M1202 359 355 227 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=108340 $D=0
M1203 360 356 228 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=112970 $D=0
M1204 231 361 359 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=108340 $D=0
M1205 232 362 360 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=112970 $D=0
M1206 361 56 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=108340 $D=0
M1207 362 56 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=112970 $D=0
M1208 161 57 363 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=108340 $D=0
M1209 162 57 364 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=112970 $D=0
M1210 365 58 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=108340 $D=0
M1211 366 58 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=112970 $D=0
M1212 367 363 217 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=108340 $D=0
M1213 368 364 218 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=112970 $D=0
M1214 161 367 723 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=108340 $D=0
M1215 162 368 724 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=112970 $D=0
M1216 369 723 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=108340 $D=0
M1217 370 724 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=112970 $D=0
M1218 367 57 369 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=108340 $D=0
M1219 368 57 370 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=112970 $D=0
M1220 369 365 227 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=108340 $D=0
M1221 370 366 228 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=112970 $D=0
M1222 231 371 369 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=108340 $D=0
M1223 232 372 370 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=112970 $D=0
M1224 371 59 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=108340 $D=0
M1225 372 59 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=112970 $D=0
M1226 161 60 373 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=108340 $D=0
M1227 162 60 374 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=112970 $D=0
M1228 375 61 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=108340 $D=0
M1229 376 61 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=112970 $D=0
M1230 377 373 217 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=108340 $D=0
M1231 378 374 218 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=112970 $D=0
M1232 161 377 725 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=108340 $D=0
M1233 162 378 726 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=112970 $D=0
M1234 379 725 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=108340 $D=0
M1235 380 726 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=112970 $D=0
M1236 377 60 379 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=108340 $D=0
M1237 378 60 380 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=112970 $D=0
M1238 379 375 227 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=108340 $D=0
M1239 380 376 228 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=112970 $D=0
M1240 231 381 379 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=108340 $D=0
M1241 232 382 380 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=112970 $D=0
M1242 381 62 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=108340 $D=0
M1243 382 62 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=112970 $D=0
M1244 161 63 383 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=108340 $D=0
M1245 162 63 384 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=112970 $D=0
M1246 385 64 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=108340 $D=0
M1247 386 64 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=112970 $D=0
M1248 387 383 217 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=108340 $D=0
M1249 388 384 218 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=112970 $D=0
M1250 161 387 727 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=108340 $D=0
M1251 162 388 728 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=112970 $D=0
M1252 389 727 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=108340 $D=0
M1253 390 728 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=112970 $D=0
M1254 387 63 389 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=108340 $D=0
M1255 388 63 390 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=112970 $D=0
M1256 389 385 227 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=108340 $D=0
M1257 390 386 228 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=112970 $D=0
M1258 231 391 389 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=108340 $D=0
M1259 232 392 390 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=112970 $D=0
M1260 391 65 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=108340 $D=0
M1261 392 65 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=112970 $D=0
M1262 161 66 393 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=108340 $D=0
M1263 162 66 394 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=112970 $D=0
M1264 395 67 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=108340 $D=0
M1265 396 67 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=112970 $D=0
M1266 397 393 217 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=108340 $D=0
M1267 398 394 218 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=112970 $D=0
M1268 161 397 729 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=108340 $D=0
M1269 162 398 730 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=112970 $D=0
M1270 399 729 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=108340 $D=0
M1271 400 730 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=112970 $D=0
M1272 397 66 399 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=108340 $D=0
M1273 398 66 400 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=112970 $D=0
M1274 399 395 227 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=108340 $D=0
M1275 400 396 228 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=112970 $D=0
M1276 231 401 399 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=108340 $D=0
M1277 232 402 400 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=112970 $D=0
M1278 401 68 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=108340 $D=0
M1279 402 68 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=112970 $D=0
M1280 161 69 403 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=108340 $D=0
M1281 162 69 404 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=112970 $D=0
M1282 405 70 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=108340 $D=0
M1283 406 70 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=112970 $D=0
M1284 407 403 217 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=108340 $D=0
M1285 408 404 218 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=112970 $D=0
M1286 161 407 731 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=108340 $D=0
M1287 162 408 732 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=112970 $D=0
M1288 409 731 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=108340 $D=0
M1289 410 732 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=112970 $D=0
M1290 407 69 409 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=108340 $D=0
M1291 408 69 410 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=112970 $D=0
M1292 409 405 227 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=108340 $D=0
M1293 410 406 228 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=112970 $D=0
M1294 231 411 409 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=108340 $D=0
M1295 232 412 410 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=112970 $D=0
M1296 411 71 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=108340 $D=0
M1297 412 71 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=112970 $D=0
M1298 161 72 413 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=108340 $D=0
M1299 162 72 414 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=112970 $D=0
M1300 415 73 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=108340 $D=0
M1301 416 73 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=112970 $D=0
M1302 417 413 217 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=108340 $D=0
M1303 418 414 218 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=112970 $D=0
M1304 161 417 733 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=108340 $D=0
M1305 162 418 734 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=112970 $D=0
M1306 419 733 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=108340 $D=0
M1307 420 734 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=112970 $D=0
M1308 417 72 419 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=108340 $D=0
M1309 418 72 420 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=112970 $D=0
M1310 419 415 227 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=108340 $D=0
M1311 420 416 228 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=112970 $D=0
M1312 231 421 419 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=108340 $D=0
M1313 232 422 420 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=112970 $D=0
M1314 421 74 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=108340 $D=0
M1315 422 74 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=112970 $D=0
M1316 161 75 423 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=108340 $D=0
M1317 162 75 424 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=112970 $D=0
M1318 425 76 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=108340 $D=0
M1319 426 76 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=112970 $D=0
M1320 427 423 217 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=108340 $D=0
M1321 428 424 218 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=112970 $D=0
M1322 161 427 735 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=108340 $D=0
M1323 162 428 736 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=112970 $D=0
M1324 429 735 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=108340 $D=0
M1325 430 736 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=112970 $D=0
M1326 427 75 429 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=108340 $D=0
M1327 428 75 430 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=112970 $D=0
M1328 429 425 227 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=108340 $D=0
M1329 430 426 228 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=112970 $D=0
M1330 231 431 429 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=108340 $D=0
M1331 232 432 430 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=112970 $D=0
M1332 431 77 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=108340 $D=0
M1333 432 77 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=112970 $D=0
M1334 161 78 433 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=108340 $D=0
M1335 162 78 434 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=112970 $D=0
M1336 435 79 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=108340 $D=0
M1337 436 79 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=112970 $D=0
M1338 437 433 217 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=108340 $D=0
M1339 438 434 218 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=112970 $D=0
M1340 161 437 737 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=108340 $D=0
M1341 162 438 738 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=112970 $D=0
M1342 439 737 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=108340 $D=0
M1343 440 738 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=112970 $D=0
M1344 437 78 439 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=108340 $D=0
M1345 438 78 440 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=112970 $D=0
M1346 439 435 227 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=108340 $D=0
M1347 440 436 228 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=112970 $D=0
M1348 231 441 439 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=108340 $D=0
M1349 232 442 440 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=112970 $D=0
M1350 441 80 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=108340 $D=0
M1351 442 80 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=112970 $D=0
M1352 161 81 443 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=108340 $D=0
M1353 162 81 444 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=112970 $D=0
M1354 445 82 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=108340 $D=0
M1355 446 82 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=112970 $D=0
M1356 447 443 217 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=108340 $D=0
M1357 448 444 218 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=112970 $D=0
M1358 161 447 739 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=108340 $D=0
M1359 162 448 740 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=112970 $D=0
M1360 449 739 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=108340 $D=0
M1361 450 740 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=112970 $D=0
M1362 447 81 449 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=108340 $D=0
M1363 448 81 450 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=112970 $D=0
M1364 449 445 227 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=108340 $D=0
M1365 450 446 228 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=112970 $D=0
M1366 231 451 449 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=108340 $D=0
M1367 232 452 450 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=112970 $D=0
M1368 451 83 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=108340 $D=0
M1369 452 83 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=112970 $D=0
M1370 161 84 453 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=108340 $D=0
M1371 162 84 454 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=112970 $D=0
M1372 455 85 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=108340 $D=0
M1373 456 85 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=112970 $D=0
M1374 457 453 217 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=108340 $D=0
M1375 458 454 218 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=112970 $D=0
M1376 161 457 741 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=108340 $D=0
M1377 162 458 742 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=112970 $D=0
M1378 459 741 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=108340 $D=0
M1379 460 742 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=112970 $D=0
M1380 457 84 459 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=108340 $D=0
M1381 458 84 460 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=112970 $D=0
M1382 459 455 227 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=108340 $D=0
M1383 460 456 228 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=112970 $D=0
M1384 231 461 459 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=108340 $D=0
M1385 232 462 460 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=112970 $D=0
M1386 461 86 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=108340 $D=0
M1387 462 86 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=112970 $D=0
M1388 161 87 463 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=108340 $D=0
M1389 162 87 464 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=112970 $D=0
M1390 465 88 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=108340 $D=0
M1391 466 88 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=112970 $D=0
M1392 467 463 217 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=108340 $D=0
M1393 468 464 218 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=112970 $D=0
M1394 161 467 743 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=108340 $D=0
M1395 162 468 744 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=112970 $D=0
M1396 469 743 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=108340 $D=0
M1397 470 744 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=112970 $D=0
M1398 467 87 469 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=108340 $D=0
M1399 468 87 470 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=112970 $D=0
M1400 469 465 227 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=108340 $D=0
M1401 470 466 228 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=112970 $D=0
M1402 231 471 469 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=108340 $D=0
M1403 232 472 470 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=112970 $D=0
M1404 471 89 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=108340 $D=0
M1405 472 89 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=112970 $D=0
M1406 161 90 473 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=108340 $D=0
M1407 162 90 474 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=112970 $D=0
M1408 475 91 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=108340 $D=0
M1409 476 91 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=112970 $D=0
M1410 477 473 217 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=108340 $D=0
M1411 478 474 218 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=112970 $D=0
M1412 161 477 745 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=108340 $D=0
M1413 162 478 746 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=112970 $D=0
M1414 479 745 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=108340 $D=0
M1415 480 746 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=112970 $D=0
M1416 477 90 479 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=108340 $D=0
M1417 478 90 480 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=112970 $D=0
M1418 479 475 227 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=108340 $D=0
M1419 480 476 228 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=112970 $D=0
M1420 231 481 479 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=108340 $D=0
M1421 232 482 480 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=112970 $D=0
M1422 481 92 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=108340 $D=0
M1423 482 92 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=112970 $D=0
M1424 161 93 483 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=108340 $D=0
M1425 162 93 484 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=112970 $D=0
M1426 485 94 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=108340 $D=0
M1427 486 94 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=112970 $D=0
M1428 487 483 217 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=108340 $D=0
M1429 488 484 218 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=112970 $D=0
M1430 161 487 747 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=108340 $D=0
M1431 162 488 748 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=112970 $D=0
M1432 489 747 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=108340 $D=0
M1433 490 748 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=112970 $D=0
M1434 487 93 489 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=108340 $D=0
M1435 488 93 490 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=112970 $D=0
M1436 489 485 227 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=108340 $D=0
M1437 490 486 228 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=112970 $D=0
M1438 231 491 489 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=108340 $D=0
M1439 232 492 490 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=112970 $D=0
M1440 491 95 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=108340 $D=0
M1441 492 95 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=112970 $D=0
M1442 161 96 493 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=108340 $D=0
M1443 162 96 494 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=112970 $D=0
M1444 495 97 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=108340 $D=0
M1445 496 97 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=112970 $D=0
M1446 497 493 217 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=108340 $D=0
M1447 498 494 218 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=112970 $D=0
M1448 161 497 749 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=108340 $D=0
M1449 162 498 750 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=112970 $D=0
M1450 499 749 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=108340 $D=0
M1451 500 750 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=112970 $D=0
M1452 497 96 499 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=108340 $D=0
M1453 498 96 500 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=112970 $D=0
M1454 499 495 227 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=108340 $D=0
M1455 500 496 228 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=112970 $D=0
M1456 231 501 499 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=108340 $D=0
M1457 232 502 500 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=112970 $D=0
M1458 501 98 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=108340 $D=0
M1459 502 98 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=112970 $D=0
M1460 161 99 503 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=108340 $D=0
M1461 162 99 504 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=112970 $D=0
M1462 505 100 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=108340 $D=0
M1463 506 100 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=112970 $D=0
M1464 507 503 217 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=108340 $D=0
M1465 508 504 218 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=112970 $D=0
M1466 161 507 751 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=108340 $D=0
M1467 162 508 752 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=112970 $D=0
M1468 509 751 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=108340 $D=0
M1469 510 752 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=112970 $D=0
M1470 507 99 509 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=108340 $D=0
M1471 508 99 510 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=112970 $D=0
M1472 509 505 227 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=108340 $D=0
M1473 510 506 228 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=112970 $D=0
M1474 231 511 509 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=108340 $D=0
M1475 232 512 510 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=112970 $D=0
M1476 511 101 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=108340 $D=0
M1477 512 101 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=112970 $D=0
M1478 161 102 513 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=108340 $D=0
M1479 162 102 514 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=112970 $D=0
M1480 515 103 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=108340 $D=0
M1481 516 103 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=112970 $D=0
M1482 517 513 217 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=108340 $D=0
M1483 518 514 218 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=112970 $D=0
M1484 161 517 753 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=108340 $D=0
M1485 162 518 754 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=112970 $D=0
M1486 519 753 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=108340 $D=0
M1487 520 754 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=112970 $D=0
M1488 517 102 519 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=108340 $D=0
M1489 518 102 520 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=112970 $D=0
M1490 519 515 227 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=108340 $D=0
M1491 520 516 228 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=112970 $D=0
M1492 231 521 519 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=108340 $D=0
M1493 232 522 520 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=112970 $D=0
M1494 521 104 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=108340 $D=0
M1495 522 104 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=112970 $D=0
M1496 161 105 523 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=108340 $D=0
M1497 162 105 524 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=112970 $D=0
M1498 525 106 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=108340 $D=0
M1499 526 106 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=112970 $D=0
M1500 527 523 217 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=108340 $D=0
M1501 528 524 218 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=112970 $D=0
M1502 161 527 755 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=108340 $D=0
M1503 162 528 756 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=112970 $D=0
M1504 529 755 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=108340 $D=0
M1505 530 756 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=112970 $D=0
M1506 527 105 529 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=108340 $D=0
M1507 528 105 530 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=112970 $D=0
M1508 529 525 227 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=108340 $D=0
M1509 530 526 228 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=112970 $D=0
M1510 231 531 529 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=108340 $D=0
M1511 232 532 530 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=112970 $D=0
M1512 531 107 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=108340 $D=0
M1513 532 107 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=112970 $D=0
M1514 161 108 533 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=108340 $D=0
M1515 162 108 534 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=112970 $D=0
M1516 535 109 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=108340 $D=0
M1517 536 109 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=112970 $D=0
M1518 4 535 227 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=108340 $D=0
M1519 8 536 228 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=112970 $D=0
M1520 231 533 4 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=108340 $D=0
M1521 232 534 8 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=112970 $D=0
M1522 161 539 537 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=108340 $D=0
M1523 162 540 538 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=112970 $D=0
M1524 539 110 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=108340 $D=0
M1525 540 110 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=112970 $D=0
M1526 757 227 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=108340 $D=0
M1527 758 228 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=112970 $D=0
M1528 541 539 757 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=108340 $D=0
M1529 542 540 758 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=112970 $D=0
M1530 161 541 543 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=108340 $D=0
M1531 162 542 544 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=112970 $D=0
M1532 759 543 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=108340 $D=0
M1533 760 544 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=112970 $D=0
M1534 541 537 759 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=108340 $D=0
M1535 542 538 760 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=112970 $D=0
M1536 161 547 545 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=108340 $D=0
M1537 162 548 546 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=112970 $D=0
M1538 547 110 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=108340 $D=0
M1539 548 110 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=112970 $D=0
M1540 761 231 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=108340 $D=0
M1541 762 232 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=112970 $D=0
M1542 549 547 761 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=108340 $D=0
M1543 550 548 762 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=112970 $D=0
M1544 161 549 111 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=108340 $D=0
M1545 162 550 112 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=112970 $D=0
M1546 763 111 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=108340 $D=0
M1547 764 112 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=112970 $D=0
M1548 549 545 763 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=108340 $D=0
M1549 550 546 764 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=112970 $D=0
M1550 551 113 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=108340 $D=0
M1551 552 113 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=112970 $D=0
M1552 553 113 543 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=108340 $D=0
M1553 554 113 544 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=112970 $D=0
M1554 114 551 553 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=108340 $D=0
M1555 115 552 554 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=112970 $D=0
M1556 555 116 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=108340 $D=0
M1557 556 116 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=112970 $D=0
M1558 557 116 111 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=108340 $D=0
M1559 558 116 112 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=112970 $D=0
M1560 765 555 557 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=108340 $D=0
M1561 766 556 558 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=112970 $D=0
M1562 161 111 765 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=108340 $D=0
M1563 162 112 766 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=112970 $D=0
M1564 559 117 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=108340 $D=0
M1565 560 117 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=112970 $D=0
M1566 561 117 557 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=108340 $D=0
M1567 562 117 558 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=112970 $D=0
M1568 9 559 561 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=108340 $D=0
M1569 10 560 562 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=112970 $D=0
M1570 564 563 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=108340 $D=0
M1571 565 118 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=112970 $D=0
M1572 161 568 566 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=108340 $D=0
M1573 162 569 567 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=112970 $D=0
M1574 570 553 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=108340 $D=0
M1575 571 554 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=112970 $D=0
M1576 568 553 563 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=108340 $D=0
M1577 569 554 118 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=112970 $D=0
M1578 564 570 568 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=108340 $D=0
M1579 565 571 569 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=112970 $D=0
M1580 572 566 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=108340 $D=0
M1581 573 567 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=112970 $D=0
M1582 574 566 561 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=108340 $D=0
M1583 563 567 562 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=112970 $D=0
M1584 553 572 574 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=108340 $D=0
M1585 554 573 563 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=112970 $D=0
M1586 575 574 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=108340 $D=0
M1587 576 563 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=112970 $D=0
M1588 577 566 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=108340 $D=0
M1589 578 567 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=112970 $D=0
M1590 579 566 575 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=108340 $D=0
M1591 580 567 576 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=112970 $D=0
M1592 561 577 579 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=108340 $D=0
M1593 562 578 580 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=112970 $D=0
M1594 788 553 161 161 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=107980 $D=0
M1595 789 554 162 162 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=112610 $D=0
M1596 581 561 788 161 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=107980 $D=0
M1597 582 562 789 162 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=112610 $D=0
M1598 583 579 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=108340 $D=0
M1599 584 580 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=112970 $D=0
M1600 585 553 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=108340 $D=0
M1601 586 554 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=112970 $D=0
M1602 161 561 585 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=108340 $D=0
M1603 162 562 586 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=112970 $D=0
M1604 587 553 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=108340 $D=0
M1605 588 554 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=112970 $D=0
M1606 161 561 587 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=108340 $D=0
M1607 162 562 588 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=112970 $D=0
M1608 790 553 161 161 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=108160 $D=0
M1609 791 554 162 162 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=112790 $D=0
M1610 591 561 790 161 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=108160 $D=0
M1611 592 562 791 162 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=112790 $D=0
M1612 161 587 591 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=108340 $D=0
M1613 162 588 592 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=112970 $D=0
M1614 593 119 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=108340 $D=0
M1615 594 119 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=112970 $D=0
M1616 595 119 581 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=108340 $D=0
M1617 596 119 582 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=112970 $D=0
M1618 585 593 595 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=108340 $D=0
M1619 586 594 596 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=112970 $D=0
M1620 597 119 583 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=108340 $D=0
M1621 598 119 584 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=112970 $D=0
M1622 591 593 597 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=108340 $D=0
M1623 592 594 598 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=112970 $D=0
M1624 599 120 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=108340 $D=0
M1625 600 120 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=112970 $D=0
M1626 601 120 597 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=108340 $D=0
M1627 602 120 598 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=112970 $D=0
M1628 595 599 601 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=108340 $D=0
M1629 596 600 602 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=112970 $D=0
M1630 11 601 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=108340 $D=0
M1631 12 602 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=112970 $D=0
M1632 603 121 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=108340 $D=0
M1633 604 121 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=112970 $D=0
M1634 605 121 122 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=108340 $D=0
M1635 606 121 123 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=112970 $D=0
M1636 124 603 605 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=108340 $D=0
M1637 125 604 606 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=112970 $D=0
M1638 607 121 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=108340 $D=0
M1639 608 121 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=112970 $D=0
M1640 613 121 127 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=108340 $D=0
M1641 614 121 129 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=112970 $D=0
M1642 130 607 613 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=108340 $D=0
M1643 128 608 614 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=112970 $D=0
M1644 615 121 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=108340 $D=0
M1645 616 121 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=112970 $D=0
M1646 133 121 131 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=108340 $D=0
M1647 133 121 132 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=112970 $D=0
M1648 134 615 133 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=108340 $D=0
M1649 135 616 133 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=112970 $D=0
M1650 617 121 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=108340 $D=0
M1651 618 121 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=112970 $D=0
M1652 619 121 136 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=108340 $D=0
M1653 620 121 8 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=112970 $D=0
M1654 137 617 619 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=108340 $D=0
M1655 138 618 620 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=112970 $D=0
M1656 621 121 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=108340 $D=0
M1657 622 121 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=112970 $D=0
M1658 623 121 4 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=108340 $D=0
M1659 624 121 8 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=112970 $D=0
M1660 139 621 623 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=108340 $D=0
M1661 140 622 624 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=112970 $D=0
M1662 161 553 778 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=108340 $D=0
M1663 162 554 779 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=112970 $D=0
M1664 125 778 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=108340 $D=0
M1665 122 779 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=112970 $D=0
M1666 625 141 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=108340 $D=0
M1667 626 141 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=112970 $D=0
M1668 143 141 125 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=108340 $D=0
M1669 144 141 122 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=112970 $D=0
M1670 605 625 143 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=108340 $D=0
M1671 606 626 144 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=112970 $D=0
M1672 627 145 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=108340 $D=0
M1673 628 145 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=112970 $D=0
M1674 126 145 143 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=108340 $D=0
M1675 146 145 144 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=112970 $D=0
M1676 613 627 126 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=108340 $D=0
M1677 614 628 146 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=112970 $D=0
M1678 629 147 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=108340 $D=0
M1679 630 147 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=112970 $D=0
M1680 142 147 126 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=108340 $D=0
M1681 148 147 146 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=112970 $D=0
M1682 133 629 142 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=108340 $D=0
M1683 133 630 148 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=112970 $D=0
M1684 631 149 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=108340 $D=0
M1685 632 149 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=112970 $D=0
M1686 150 149 142 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=108340 $D=0
M1687 151 149 148 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=112970 $D=0
M1688 619 631 150 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=108340 $D=0
M1689 620 632 151 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=112970 $D=0
M1690 633 152 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=108340 $D=0
M1691 634 152 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=112970 $D=0
M1692 203 152 150 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=108340 $D=0
M1693 204 152 151 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=112970 $D=0
M1694 623 633 203 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=108340 $D=0
M1695 624 634 204 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=112970 $D=0
M1696 635 153 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=108340 $D=0
M1697 636 153 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=112970 $D=0
M1698 637 153 111 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=108340 $D=0
M1699 638 153 112 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=112970 $D=0
M1700 9 635 637 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=108340 $D=0
M1701 10 636 638 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=112970 $D=0
M1702 639 543 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=108340 $D=0
M1703 640 544 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=112970 $D=0
M1704 161 637 639 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=108340 $D=0
M1705 162 638 640 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=112970 $D=0
M1706 792 543 161 161 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=108160 $D=0
M1707 793 544 162 162 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=112790 $D=0
M1708 643 637 792 161 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=108160 $D=0
M1709 644 638 793 162 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=112790 $D=0
M1710 161 639 643 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=108340 $D=0
M1711 162 640 644 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=112970 $D=0
M1712 780 645 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=108340 $D=0
M1713 781 646 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=112970 $D=0
M1714 161 643 780 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=108340 $D=0
M1715 162 644 781 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=112970 $D=0
M1716 646 780 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=108340 $D=0
M1717 154 781 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=112970 $D=0
M1718 794 543 161 161 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=107980 $D=0
M1719 795 544 162 162 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=112610 $D=0
M1720 647 649 794 161 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=107980 $D=0
M1721 648 650 795 162 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=112610 $D=0
M1722 649 637 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=108340 $D=0
M1723 650 638 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=112970 $D=0
M1724 651 647 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=108340 $D=0
M1725 652 648 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=112970 $D=0
M1726 161 645 651 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=108340 $D=0
M1727 162 646 652 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=112970 $D=0
M1728 654 155 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=108340 $D=0
M1729 655 653 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=112970 $D=0
M1730 653 651 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=108340 $D=0
M1731 156 652 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=112970 $D=0
M1732 161 654 653 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=108340 $D=0
M1733 162 655 156 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=112970 $D=0
M1734 657 656 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=108340 $D=0
M1735 658 157 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=112970 $D=0
M1736 161 661 659 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=108340 $D=0
M1737 162 662 660 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=112970 $D=0
M1738 663 114 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=108340 $D=0
M1739 664 115 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=112970 $D=0
M1740 661 114 656 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=108340 $D=0
M1741 662 115 157 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=112970 $D=0
M1742 657 663 661 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=108340 $D=0
M1743 658 664 662 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=112970 $D=0
M1744 665 659 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=108340 $D=0
M1745 666 660 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=112970 $D=0
M1746 158 659 4 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=108340 $D=0
M1747 656 660 8 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=112970 $D=0
M1748 114 665 158 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=108340 $D=0
M1749 115 666 656 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=112970 $D=0
M1750 667 158 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=108340 $D=0
M1751 668 656 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=112970 $D=0
M1752 669 659 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=108340 $D=0
M1753 670 660 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=112970 $D=0
M1754 205 659 667 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=108340 $D=0
M1755 206 660 668 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=112970 $D=0
M1756 4 669 205 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=108340 $D=0
M1757 8 670 206 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=112970 $D=0
M1758 671 159 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=108340 $D=0
M1759 672 159 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=112970 $D=0
M1760 673 159 205 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=108340 $D=0
M1761 674 159 206 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=112970 $D=0
M1762 11 671 673 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=108340 $D=0
M1763 12 672 674 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=112970 $D=0
M1764 675 160 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=108340 $D=0
M1765 676 160 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=112970 $D=0
M1766 160 160 673 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=108340 $D=0
M1767 160 160 674 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=112970 $D=0
M1768 4 675 160 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=108340 $D=0
M1769 8 676 160 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=112970 $D=0
M1770 677 110 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=108340 $D=0
M1771 678 110 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=112970 $D=0
M1772 161 677 679 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=108340 $D=0
M1773 162 678 680 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=112970 $D=0
M1774 681 110 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=108340 $D=0
M1775 682 110 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=112970 $D=0
M1776 683 679 160 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=108340 $D=0
M1777 684 680 160 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=112970 $D=0
M1778 161 683 782 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=108340 $D=0
M1779 162 684 783 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=112970 $D=0
M1780 685 782 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=108340 $D=0
M1781 686 783 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=112970 $D=0
M1782 683 677 685 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=108340 $D=0
M1783 684 678 686 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=112970 $D=0
M1784 687 681 685 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=108340 $D=0
M1785 688 682 686 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=112970 $D=0
M1786 161 691 689 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=108340 $D=0
M1787 162 692 690 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=112970 $D=0
M1788 691 110 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=108340 $D=0
M1789 692 110 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=112970 $D=0
M1790 784 687 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=108340 $D=0
M1791 785 688 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=112970 $D=0
M1792 693 691 784 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=108340 $D=0
M1793 694 692 785 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=112970 $D=0
M1794 161 693 114 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=108340 $D=0
M1795 162 694 115 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=112970 $D=0
M1796 786 114 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=108340 $D=0
M1797 787 115 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=112970 $D=0
M1798 693 689 786 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=108340 $D=0
M1799 694 690 787 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=112970 $D=0
.ENDS
***************************************
.SUBCKT ICV_28 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164
** N=806 EP=164 IP=1514 FDC=1800
M0 177 1 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=97830 $D=1
M1 178 1 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=102460 $D=1
M2 179 177 2 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=97830 $D=1
M3 180 178 3 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=102460 $D=1
M4 5 1 179 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=97830 $D=1
M5 6 1 180 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=102460 $D=1
M6 181 177 4 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=97830 $D=1
M7 182 178 4 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=102460 $D=1
M8 2 1 181 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=97830 $D=1
M9 3 1 182 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=102460 $D=1
M10 183 177 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=97830 $D=1
M11 184 178 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=102460 $D=1
M12 2 1 183 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=97830 $D=1
M13 3 1 184 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=102460 $D=1
M14 187 185 183 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=97830 $D=1
M15 188 186 184 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=102460 $D=1
M16 185 7 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=97830 $D=1
M17 186 7 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=102460 $D=1
M18 189 185 181 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=97830 $D=1
M19 190 186 182 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=102460 $D=1
M20 179 7 189 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=97830 $D=1
M21 180 7 190 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=102460 $D=1
M22 191 8 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=97830 $D=1
M23 192 8 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=102460 $D=1
M24 193 191 189 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=97830 $D=1
M25 194 192 190 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=102460 $D=1
M26 187 8 193 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=97830 $D=1
M27 188 8 194 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=102460 $D=1
M28 195 9 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=97830 $D=1
M29 196 9 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=102460 $D=1
M30 197 195 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=97830 $D=1
M31 198 196 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=102460 $D=1
M32 10 9 197 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=97830 $D=1
M33 11 9 198 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=102460 $D=1
M34 199 195 12 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=97830 $D=1
M35 200 196 13 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=102460 $D=1
M36 201 9 199 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=97830 $D=1
M37 202 9 200 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=102460 $D=1
M38 205 195 203 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=97830 $D=1
M39 206 196 204 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=102460 $D=1
M40 193 9 205 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=97830 $D=1
M41 194 9 206 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=102460 $D=1
M42 209 207 205 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=97830 $D=1
M43 210 208 206 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=102460 $D=1
M44 207 14 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=97830 $D=1
M45 208 14 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=102460 $D=1
M46 211 207 199 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=97830 $D=1
M47 212 208 200 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=102460 $D=1
M48 197 14 211 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=97830 $D=1
M49 198 14 212 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=102460 $D=1
M50 213 15 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=97830 $D=1
M51 214 15 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=102460 $D=1
M52 215 213 211 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=97830 $D=1
M53 216 214 212 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=102460 $D=1
M54 209 15 215 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=97830 $D=1
M55 210 15 216 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=102460 $D=1
M56 5 16 217 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=97830 $D=1
M57 6 16 218 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=102460 $D=1
M58 219 17 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=97830 $D=1
M59 220 17 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=102460 $D=1
M60 221 16 215 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=97830 $D=1
M61 222 16 216 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=102460 $D=1
M62 5 221 693 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=97830 $D=1
M63 6 222 694 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=102460 $D=1
M64 223 693 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=97830 $D=1
M65 224 694 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=102460 $D=1
M66 221 217 223 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=97830 $D=1
M67 222 218 224 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=102460 $D=1
M68 223 17 225 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=97830 $D=1
M69 224 17 226 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=102460 $D=1
M70 229 18 223 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=97830 $D=1
M71 230 18 224 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=102460 $D=1
M72 227 18 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=97830 $D=1
M73 228 18 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=102460 $D=1
M74 5 19 231 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=97830 $D=1
M75 6 19 232 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=102460 $D=1
M76 233 20 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=97830 $D=1
M77 234 20 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=102460 $D=1
M78 235 19 215 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=97830 $D=1
M79 236 19 216 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=102460 $D=1
M80 5 235 695 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=97830 $D=1
M81 6 236 696 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=102460 $D=1
M82 237 695 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=97830 $D=1
M83 238 696 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=102460 $D=1
M84 235 231 237 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=97830 $D=1
M85 236 232 238 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=102460 $D=1
M86 237 20 225 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=97830 $D=1
M87 238 20 226 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=102460 $D=1
M88 229 21 237 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=97830 $D=1
M89 230 21 238 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=102460 $D=1
M90 239 21 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=97830 $D=1
M91 240 21 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=102460 $D=1
M92 5 22 241 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=97830 $D=1
M93 6 22 242 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=102460 $D=1
M94 243 23 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=97830 $D=1
M95 244 23 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=102460 $D=1
M96 245 22 215 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=97830 $D=1
M97 246 22 216 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=102460 $D=1
M98 5 245 697 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=97830 $D=1
M99 6 246 698 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=102460 $D=1
M100 247 697 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=97830 $D=1
M101 248 698 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=102460 $D=1
M102 245 241 247 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=97830 $D=1
M103 246 242 248 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=102460 $D=1
M104 247 23 225 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=97830 $D=1
M105 248 23 226 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=102460 $D=1
M106 229 24 247 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=97830 $D=1
M107 230 24 248 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=102460 $D=1
M108 249 24 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=97830 $D=1
M109 250 24 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=102460 $D=1
M110 5 25 251 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=97830 $D=1
M111 6 25 252 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=102460 $D=1
M112 253 26 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=97830 $D=1
M113 254 26 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=102460 $D=1
M114 255 25 215 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=97830 $D=1
M115 256 25 216 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=102460 $D=1
M116 5 255 699 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=97830 $D=1
M117 6 256 700 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=102460 $D=1
M118 257 699 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=97830 $D=1
M119 258 700 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=102460 $D=1
M120 255 251 257 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=97830 $D=1
M121 256 252 258 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=102460 $D=1
M122 257 26 225 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=97830 $D=1
M123 258 26 226 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=102460 $D=1
M124 229 27 257 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=97830 $D=1
M125 230 27 258 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=102460 $D=1
M126 259 27 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=97830 $D=1
M127 260 27 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=102460 $D=1
M128 5 28 261 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=97830 $D=1
M129 6 28 262 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=102460 $D=1
M130 263 29 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=97830 $D=1
M131 264 29 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=102460 $D=1
M132 265 28 215 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=97830 $D=1
M133 266 28 216 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=102460 $D=1
M134 5 265 701 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=97830 $D=1
M135 6 266 702 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=102460 $D=1
M136 267 701 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=97830 $D=1
M137 268 702 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=102460 $D=1
M138 265 261 267 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=97830 $D=1
M139 266 262 268 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=102460 $D=1
M140 267 29 225 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=97830 $D=1
M141 268 29 226 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=102460 $D=1
M142 229 30 267 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=97830 $D=1
M143 230 30 268 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=102460 $D=1
M144 269 30 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=97830 $D=1
M145 270 30 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=102460 $D=1
M146 5 31 271 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=97830 $D=1
M147 6 31 272 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=102460 $D=1
M148 273 32 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=97830 $D=1
M149 274 32 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=102460 $D=1
M150 275 31 215 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=97830 $D=1
M151 276 31 216 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=102460 $D=1
M152 5 275 703 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=97830 $D=1
M153 6 276 704 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=102460 $D=1
M154 277 703 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=97830 $D=1
M155 278 704 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=102460 $D=1
M156 275 271 277 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=97830 $D=1
M157 276 272 278 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=102460 $D=1
M158 277 32 225 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=97830 $D=1
M159 278 32 226 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=102460 $D=1
M160 229 33 277 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=97830 $D=1
M161 230 33 278 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=102460 $D=1
M162 279 33 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=97830 $D=1
M163 280 33 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=102460 $D=1
M164 5 34 281 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=97830 $D=1
M165 6 34 282 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=102460 $D=1
M166 283 35 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=97830 $D=1
M167 284 35 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=102460 $D=1
M168 285 34 215 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=97830 $D=1
M169 286 34 216 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=102460 $D=1
M170 5 285 705 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=97830 $D=1
M171 6 286 706 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=102460 $D=1
M172 287 705 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=97830 $D=1
M173 288 706 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=102460 $D=1
M174 285 281 287 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=97830 $D=1
M175 286 282 288 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=102460 $D=1
M176 287 35 225 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=97830 $D=1
M177 288 35 226 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=102460 $D=1
M178 229 36 287 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=97830 $D=1
M179 230 36 288 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=102460 $D=1
M180 289 36 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=97830 $D=1
M181 290 36 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=102460 $D=1
M182 5 37 291 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=97830 $D=1
M183 6 37 292 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=102460 $D=1
M184 293 38 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=97830 $D=1
M185 294 38 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=102460 $D=1
M186 295 37 215 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=97830 $D=1
M187 296 37 216 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=102460 $D=1
M188 5 295 707 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=97830 $D=1
M189 6 296 708 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=102460 $D=1
M190 297 707 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=97830 $D=1
M191 298 708 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=102460 $D=1
M192 295 291 297 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=97830 $D=1
M193 296 292 298 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=102460 $D=1
M194 297 38 225 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=97830 $D=1
M195 298 38 226 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=102460 $D=1
M196 229 39 297 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=97830 $D=1
M197 230 39 298 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=102460 $D=1
M198 299 39 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=97830 $D=1
M199 300 39 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=102460 $D=1
M200 5 40 301 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=97830 $D=1
M201 6 40 302 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=102460 $D=1
M202 303 41 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=97830 $D=1
M203 304 41 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=102460 $D=1
M204 305 40 215 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=97830 $D=1
M205 306 40 216 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=102460 $D=1
M206 5 305 709 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=97830 $D=1
M207 6 306 710 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=102460 $D=1
M208 307 709 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=97830 $D=1
M209 308 710 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=102460 $D=1
M210 305 301 307 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=97830 $D=1
M211 306 302 308 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=102460 $D=1
M212 307 41 225 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=97830 $D=1
M213 308 41 226 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=102460 $D=1
M214 229 42 307 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=97830 $D=1
M215 230 42 308 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=102460 $D=1
M216 309 42 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=97830 $D=1
M217 310 42 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=102460 $D=1
M218 5 43 311 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=97830 $D=1
M219 6 43 312 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=102460 $D=1
M220 313 44 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=97830 $D=1
M221 314 44 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=102460 $D=1
M222 315 43 215 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=97830 $D=1
M223 316 43 216 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=102460 $D=1
M224 5 315 711 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=97830 $D=1
M225 6 316 712 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=102460 $D=1
M226 317 711 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=97830 $D=1
M227 318 712 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=102460 $D=1
M228 315 311 317 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=97830 $D=1
M229 316 312 318 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=102460 $D=1
M230 317 44 225 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=97830 $D=1
M231 318 44 226 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=102460 $D=1
M232 229 45 317 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=97830 $D=1
M233 230 45 318 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=102460 $D=1
M234 319 45 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=97830 $D=1
M235 320 45 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=102460 $D=1
M236 5 46 321 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=97830 $D=1
M237 6 46 322 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=102460 $D=1
M238 323 47 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=97830 $D=1
M239 324 47 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=102460 $D=1
M240 325 46 215 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=97830 $D=1
M241 326 46 216 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=102460 $D=1
M242 5 325 713 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=97830 $D=1
M243 6 326 714 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=102460 $D=1
M244 327 713 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=97830 $D=1
M245 328 714 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=102460 $D=1
M246 325 321 327 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=97830 $D=1
M247 326 322 328 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=102460 $D=1
M248 327 47 225 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=97830 $D=1
M249 328 47 226 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=102460 $D=1
M250 229 48 327 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=97830 $D=1
M251 230 48 328 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=102460 $D=1
M252 329 48 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=97830 $D=1
M253 330 48 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=102460 $D=1
M254 5 49 331 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=97830 $D=1
M255 6 49 332 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=102460 $D=1
M256 333 50 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=97830 $D=1
M257 334 50 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=102460 $D=1
M258 335 49 215 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=97830 $D=1
M259 336 49 216 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=102460 $D=1
M260 5 335 715 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=97830 $D=1
M261 6 336 716 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=102460 $D=1
M262 337 715 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=97830 $D=1
M263 338 716 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=102460 $D=1
M264 335 331 337 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=97830 $D=1
M265 336 332 338 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=102460 $D=1
M266 337 50 225 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=97830 $D=1
M267 338 50 226 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=102460 $D=1
M268 229 51 337 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=97830 $D=1
M269 230 51 338 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=102460 $D=1
M270 339 51 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=97830 $D=1
M271 340 51 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=102460 $D=1
M272 5 52 341 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=97830 $D=1
M273 6 52 342 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=102460 $D=1
M274 343 53 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=97830 $D=1
M275 344 53 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=102460 $D=1
M276 345 52 215 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=97830 $D=1
M277 346 52 216 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=102460 $D=1
M278 5 345 717 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=97830 $D=1
M279 6 346 718 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=102460 $D=1
M280 347 717 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=97830 $D=1
M281 348 718 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=102460 $D=1
M282 345 341 347 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=97830 $D=1
M283 346 342 348 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=102460 $D=1
M284 347 53 225 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=97830 $D=1
M285 348 53 226 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=102460 $D=1
M286 229 54 347 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=97830 $D=1
M287 230 54 348 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=102460 $D=1
M288 349 54 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=97830 $D=1
M289 350 54 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=102460 $D=1
M290 5 55 351 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=97830 $D=1
M291 6 55 352 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=102460 $D=1
M292 353 56 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=97830 $D=1
M293 354 56 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=102460 $D=1
M294 355 55 215 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=97830 $D=1
M295 356 55 216 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=102460 $D=1
M296 5 355 719 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=97830 $D=1
M297 6 356 720 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=102460 $D=1
M298 357 719 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=97830 $D=1
M299 358 720 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=102460 $D=1
M300 355 351 357 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=97830 $D=1
M301 356 352 358 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=102460 $D=1
M302 357 56 225 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=97830 $D=1
M303 358 56 226 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=102460 $D=1
M304 229 57 357 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=97830 $D=1
M305 230 57 358 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=102460 $D=1
M306 359 57 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=97830 $D=1
M307 360 57 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=102460 $D=1
M308 5 58 361 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=97830 $D=1
M309 6 58 362 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=102460 $D=1
M310 363 59 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=97830 $D=1
M311 364 59 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=102460 $D=1
M312 365 58 215 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=97830 $D=1
M313 366 58 216 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=102460 $D=1
M314 5 365 721 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=97830 $D=1
M315 6 366 722 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=102460 $D=1
M316 367 721 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=97830 $D=1
M317 368 722 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=102460 $D=1
M318 365 361 367 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=97830 $D=1
M319 366 362 368 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=102460 $D=1
M320 367 59 225 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=97830 $D=1
M321 368 59 226 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=102460 $D=1
M322 229 60 367 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=97830 $D=1
M323 230 60 368 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=102460 $D=1
M324 369 60 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=97830 $D=1
M325 370 60 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=102460 $D=1
M326 5 61 371 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=97830 $D=1
M327 6 61 372 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=102460 $D=1
M328 373 62 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=97830 $D=1
M329 374 62 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=102460 $D=1
M330 375 61 215 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=97830 $D=1
M331 376 61 216 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=102460 $D=1
M332 5 375 723 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=97830 $D=1
M333 6 376 724 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=102460 $D=1
M334 377 723 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=97830 $D=1
M335 378 724 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=102460 $D=1
M336 375 371 377 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=97830 $D=1
M337 376 372 378 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=102460 $D=1
M338 377 62 225 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=97830 $D=1
M339 378 62 226 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=102460 $D=1
M340 229 63 377 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=97830 $D=1
M341 230 63 378 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=102460 $D=1
M342 379 63 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=97830 $D=1
M343 380 63 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=102460 $D=1
M344 5 64 381 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=97830 $D=1
M345 6 64 382 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=102460 $D=1
M346 383 65 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=97830 $D=1
M347 384 65 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=102460 $D=1
M348 385 64 215 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=97830 $D=1
M349 386 64 216 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=102460 $D=1
M350 5 385 725 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=97830 $D=1
M351 6 386 726 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=102460 $D=1
M352 387 725 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=97830 $D=1
M353 388 726 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=102460 $D=1
M354 385 381 387 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=97830 $D=1
M355 386 382 388 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=102460 $D=1
M356 387 65 225 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=97830 $D=1
M357 388 65 226 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=102460 $D=1
M358 229 66 387 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=97830 $D=1
M359 230 66 388 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=102460 $D=1
M360 389 66 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=97830 $D=1
M361 390 66 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=102460 $D=1
M362 5 67 391 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=97830 $D=1
M363 6 67 392 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=102460 $D=1
M364 393 68 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=97830 $D=1
M365 394 68 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=102460 $D=1
M366 395 67 215 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=97830 $D=1
M367 396 67 216 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=102460 $D=1
M368 5 395 727 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=97830 $D=1
M369 6 396 728 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=102460 $D=1
M370 397 727 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=97830 $D=1
M371 398 728 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=102460 $D=1
M372 395 391 397 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=97830 $D=1
M373 396 392 398 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=102460 $D=1
M374 397 68 225 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=97830 $D=1
M375 398 68 226 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=102460 $D=1
M376 229 69 397 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=97830 $D=1
M377 230 69 398 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=102460 $D=1
M378 399 69 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=97830 $D=1
M379 400 69 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=102460 $D=1
M380 5 70 401 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=97830 $D=1
M381 6 70 402 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=102460 $D=1
M382 403 71 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=97830 $D=1
M383 404 71 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=102460 $D=1
M384 405 70 215 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=97830 $D=1
M385 406 70 216 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=102460 $D=1
M386 5 405 729 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=97830 $D=1
M387 6 406 730 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=102460 $D=1
M388 407 729 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=97830 $D=1
M389 408 730 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=102460 $D=1
M390 405 401 407 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=97830 $D=1
M391 406 402 408 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=102460 $D=1
M392 407 71 225 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=97830 $D=1
M393 408 71 226 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=102460 $D=1
M394 229 72 407 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=97830 $D=1
M395 230 72 408 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=102460 $D=1
M396 409 72 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=97830 $D=1
M397 410 72 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=102460 $D=1
M398 5 73 411 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=97830 $D=1
M399 6 73 412 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=102460 $D=1
M400 413 74 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=97830 $D=1
M401 414 74 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=102460 $D=1
M402 415 73 215 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=97830 $D=1
M403 416 73 216 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=102460 $D=1
M404 5 415 731 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=97830 $D=1
M405 6 416 732 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=102460 $D=1
M406 417 731 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=97830 $D=1
M407 418 732 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=102460 $D=1
M408 415 411 417 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=97830 $D=1
M409 416 412 418 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=102460 $D=1
M410 417 74 225 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=97830 $D=1
M411 418 74 226 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=102460 $D=1
M412 229 75 417 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=97830 $D=1
M413 230 75 418 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=102460 $D=1
M414 419 75 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=97830 $D=1
M415 420 75 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=102460 $D=1
M416 5 76 421 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=97830 $D=1
M417 6 76 422 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=102460 $D=1
M418 423 77 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=97830 $D=1
M419 424 77 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=102460 $D=1
M420 425 76 215 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=97830 $D=1
M421 426 76 216 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=102460 $D=1
M422 5 425 733 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=97830 $D=1
M423 6 426 734 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=102460 $D=1
M424 427 733 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=97830 $D=1
M425 428 734 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=102460 $D=1
M426 425 421 427 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=97830 $D=1
M427 426 422 428 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=102460 $D=1
M428 427 77 225 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=97830 $D=1
M429 428 77 226 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=102460 $D=1
M430 229 78 427 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=97830 $D=1
M431 230 78 428 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=102460 $D=1
M432 429 78 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=97830 $D=1
M433 430 78 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=102460 $D=1
M434 5 79 431 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=97830 $D=1
M435 6 79 432 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=102460 $D=1
M436 433 80 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=97830 $D=1
M437 434 80 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=102460 $D=1
M438 435 79 215 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=97830 $D=1
M439 436 79 216 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=102460 $D=1
M440 5 435 735 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=97830 $D=1
M441 6 436 736 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=102460 $D=1
M442 437 735 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=97830 $D=1
M443 438 736 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=102460 $D=1
M444 435 431 437 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=97830 $D=1
M445 436 432 438 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=102460 $D=1
M446 437 80 225 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=97830 $D=1
M447 438 80 226 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=102460 $D=1
M448 229 81 437 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=97830 $D=1
M449 230 81 438 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=102460 $D=1
M450 439 81 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=97830 $D=1
M451 440 81 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=102460 $D=1
M452 5 82 441 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=97830 $D=1
M453 6 82 442 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=102460 $D=1
M454 443 83 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=97830 $D=1
M455 444 83 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=102460 $D=1
M456 445 82 215 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=97830 $D=1
M457 446 82 216 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=102460 $D=1
M458 5 445 737 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=97830 $D=1
M459 6 446 738 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=102460 $D=1
M460 447 737 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=97830 $D=1
M461 448 738 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=102460 $D=1
M462 445 441 447 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=97830 $D=1
M463 446 442 448 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=102460 $D=1
M464 447 83 225 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=97830 $D=1
M465 448 83 226 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=102460 $D=1
M466 229 84 447 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=97830 $D=1
M467 230 84 448 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=102460 $D=1
M468 449 84 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=97830 $D=1
M469 450 84 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=102460 $D=1
M470 5 85 451 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=97830 $D=1
M471 6 85 452 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=102460 $D=1
M472 453 86 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=97830 $D=1
M473 454 86 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=102460 $D=1
M474 455 85 215 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=97830 $D=1
M475 456 85 216 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=102460 $D=1
M476 5 455 739 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=97830 $D=1
M477 6 456 740 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=102460 $D=1
M478 457 739 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=97830 $D=1
M479 458 740 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=102460 $D=1
M480 455 451 457 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=97830 $D=1
M481 456 452 458 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=102460 $D=1
M482 457 86 225 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=97830 $D=1
M483 458 86 226 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=102460 $D=1
M484 229 87 457 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=97830 $D=1
M485 230 87 458 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=102460 $D=1
M486 459 87 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=97830 $D=1
M487 460 87 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=102460 $D=1
M488 5 88 461 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=97830 $D=1
M489 6 88 462 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=102460 $D=1
M490 463 89 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=97830 $D=1
M491 464 89 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=102460 $D=1
M492 465 88 215 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=97830 $D=1
M493 466 88 216 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=102460 $D=1
M494 5 465 741 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=97830 $D=1
M495 6 466 742 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=102460 $D=1
M496 467 741 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=97830 $D=1
M497 468 742 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=102460 $D=1
M498 465 461 467 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=97830 $D=1
M499 466 462 468 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=102460 $D=1
M500 467 89 225 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=97830 $D=1
M501 468 89 226 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=102460 $D=1
M502 229 90 467 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=97830 $D=1
M503 230 90 468 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=102460 $D=1
M504 469 90 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=97830 $D=1
M505 470 90 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=102460 $D=1
M506 5 91 471 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=97830 $D=1
M507 6 91 472 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=102460 $D=1
M508 473 92 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=97830 $D=1
M509 474 92 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=102460 $D=1
M510 475 91 215 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=97830 $D=1
M511 476 91 216 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=102460 $D=1
M512 5 475 743 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=97830 $D=1
M513 6 476 744 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=102460 $D=1
M514 477 743 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=97830 $D=1
M515 478 744 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=102460 $D=1
M516 475 471 477 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=97830 $D=1
M517 476 472 478 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=102460 $D=1
M518 477 92 225 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=97830 $D=1
M519 478 92 226 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=102460 $D=1
M520 229 93 477 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=97830 $D=1
M521 230 93 478 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=102460 $D=1
M522 479 93 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=97830 $D=1
M523 480 93 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=102460 $D=1
M524 5 94 481 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=97830 $D=1
M525 6 94 482 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=102460 $D=1
M526 483 95 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=97830 $D=1
M527 484 95 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=102460 $D=1
M528 485 94 215 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=97830 $D=1
M529 486 94 216 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=102460 $D=1
M530 5 485 745 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=97830 $D=1
M531 6 486 746 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=102460 $D=1
M532 487 745 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=97830 $D=1
M533 488 746 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=102460 $D=1
M534 485 481 487 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=97830 $D=1
M535 486 482 488 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=102460 $D=1
M536 487 95 225 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=97830 $D=1
M537 488 95 226 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=102460 $D=1
M538 229 96 487 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=97830 $D=1
M539 230 96 488 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=102460 $D=1
M540 489 96 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=97830 $D=1
M541 490 96 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=102460 $D=1
M542 5 97 491 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=97830 $D=1
M543 6 97 492 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=102460 $D=1
M544 493 98 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=97830 $D=1
M545 494 98 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=102460 $D=1
M546 495 97 215 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=97830 $D=1
M547 496 97 216 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=102460 $D=1
M548 5 495 747 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=97830 $D=1
M549 6 496 748 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=102460 $D=1
M550 497 747 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=97830 $D=1
M551 498 748 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=102460 $D=1
M552 495 491 497 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=97830 $D=1
M553 496 492 498 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=102460 $D=1
M554 497 98 225 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=97830 $D=1
M555 498 98 226 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=102460 $D=1
M556 229 99 497 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=97830 $D=1
M557 230 99 498 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=102460 $D=1
M558 499 99 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=97830 $D=1
M559 500 99 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=102460 $D=1
M560 5 100 501 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=97830 $D=1
M561 6 100 502 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=102460 $D=1
M562 503 101 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=97830 $D=1
M563 504 101 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=102460 $D=1
M564 505 100 215 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=97830 $D=1
M565 506 100 216 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=102460 $D=1
M566 5 505 749 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=97830 $D=1
M567 6 506 750 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=102460 $D=1
M568 507 749 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=97830 $D=1
M569 508 750 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=102460 $D=1
M570 505 501 507 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=97830 $D=1
M571 506 502 508 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=102460 $D=1
M572 507 101 225 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=97830 $D=1
M573 508 101 226 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=102460 $D=1
M574 229 102 507 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=97830 $D=1
M575 230 102 508 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=102460 $D=1
M576 509 102 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=97830 $D=1
M577 510 102 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=102460 $D=1
M578 5 103 511 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=97830 $D=1
M579 6 103 512 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=102460 $D=1
M580 513 104 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=97830 $D=1
M581 514 104 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=102460 $D=1
M582 515 103 215 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=97830 $D=1
M583 516 103 216 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=102460 $D=1
M584 5 515 751 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=97830 $D=1
M585 6 516 752 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=102460 $D=1
M586 517 751 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=97830 $D=1
M587 518 752 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=102460 $D=1
M588 515 511 517 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=97830 $D=1
M589 516 512 518 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=102460 $D=1
M590 517 104 225 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=97830 $D=1
M591 518 104 226 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=102460 $D=1
M592 229 105 517 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=97830 $D=1
M593 230 105 518 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=102460 $D=1
M594 519 105 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=97830 $D=1
M595 520 105 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=102460 $D=1
M596 5 106 521 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=97830 $D=1
M597 6 106 522 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=102460 $D=1
M598 523 107 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=97830 $D=1
M599 524 107 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=102460 $D=1
M600 525 106 215 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=97830 $D=1
M601 526 106 216 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=102460 $D=1
M602 5 525 753 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=97830 $D=1
M603 6 526 754 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=102460 $D=1
M604 527 753 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=97830 $D=1
M605 528 754 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=102460 $D=1
M606 525 521 527 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=97830 $D=1
M607 526 522 528 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=102460 $D=1
M608 527 107 225 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=97830 $D=1
M609 528 107 226 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=102460 $D=1
M610 229 108 527 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=97830 $D=1
M611 230 108 528 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=102460 $D=1
M612 529 108 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=97830 $D=1
M613 530 108 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=102460 $D=1
M614 5 109 531 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=97830 $D=1
M615 6 109 532 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=102460 $D=1
M616 533 110 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=97830 $D=1
M617 534 110 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=102460 $D=1
M618 5 110 225 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=97830 $D=1
M619 6 110 226 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=102460 $D=1
M620 229 109 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=97830 $D=1
M621 230 109 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=102460 $D=1
M622 5 537 535 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=97830 $D=1
M623 6 538 536 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=102460 $D=1
M624 537 111 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=97830 $D=1
M625 538 111 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=102460 $D=1
M626 755 225 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=97830 $D=1
M627 756 226 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=102460 $D=1
M628 539 535 755 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=97830 $D=1
M629 540 536 756 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=102460 $D=1
M630 5 539 541 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=97830 $D=1
M631 6 540 542 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=102460 $D=1
M632 757 541 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=97830 $D=1
M633 758 542 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=102460 $D=1
M634 539 537 757 5 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=97830 $D=1
M635 540 538 758 6 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=102460 $D=1
M636 5 545 543 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=97830 $D=1
M637 6 546 544 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=102460 $D=1
M638 545 111 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=97830 $D=1
M639 546 111 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=102460 $D=1
M640 759 229 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=97830 $D=1
M641 760 230 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=102460 $D=1
M642 547 543 759 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=97830 $D=1
M643 548 544 760 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=102460 $D=1
M644 5 547 112 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=97830 $D=1
M645 6 548 113 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=102460 $D=1
M646 761 112 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=97830 $D=1
M647 762 113 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=102460 $D=1
M648 547 545 761 5 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=97830 $D=1
M649 548 546 762 6 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=102460 $D=1
M650 549 114 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=97830 $D=1
M651 550 114 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=102460 $D=1
M652 551 549 541 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=97830 $D=1
M653 552 550 542 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=102460 $D=1
M654 115 114 551 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=97830 $D=1
M655 116 114 552 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=102460 $D=1
M656 553 117 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=97830 $D=1
M657 554 117 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=102460 $D=1
M658 555 553 112 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=97830 $D=1
M659 556 554 113 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=102460 $D=1
M660 763 117 555 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=97830 $D=1
M661 764 117 556 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=102460 $D=1
M662 5 112 763 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=97830 $D=1
M663 6 113 764 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=102460 $D=1
M664 557 118 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=97830 $D=1
M665 558 118 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=102460 $D=1
M666 559 557 555 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=97830 $D=1
M667 560 558 556 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=102460 $D=1
M668 10 118 559 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=97830 $D=1
M669 11 118 560 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=102460 $D=1
M670 562 561 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=97830 $D=1
M671 563 119 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=102460 $D=1
M672 5 566 564 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=97830 $D=1
M673 6 567 565 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=102460 $D=1
M674 568 551 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=97830 $D=1
M675 569 552 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=102460 $D=1
M676 566 568 561 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=97830 $D=1
M677 567 569 119 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=102460 $D=1
M678 562 551 566 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=97830 $D=1
M679 563 552 567 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=102460 $D=1
M680 570 564 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=97830 $D=1
M681 571 565 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=102460 $D=1
M682 120 570 559 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=97830 $D=1
M683 561 571 560 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=102460 $D=1
M684 551 564 120 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=97830 $D=1
M685 552 565 561 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=102460 $D=1
M686 572 120 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=97830 $D=1
M687 573 561 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=102460 $D=1
M688 574 564 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=97830 $D=1
M689 575 565 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=102460 $D=1
M690 576 574 572 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=97830 $D=1
M691 577 575 573 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=102460 $D=1
M692 559 564 576 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=97830 $D=1
M693 560 565 577 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=102460 $D=1
M694 578 551 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=97830 $D=1
M695 579 552 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=102460 $D=1
M696 5 559 578 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=97830 $D=1
M697 6 560 579 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=102460 $D=1
M698 580 576 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=97830 $D=1
M699 581 577 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=102460 $D=1
M700 795 551 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=97830 $D=1
M701 796 552 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=102460 $D=1
M702 582 559 795 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=97830 $D=1
M703 583 560 796 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=102460 $D=1
M704 797 551 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=97830 $D=1
M705 798 552 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=102460 $D=1
M706 584 559 797 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=97830 $D=1
M707 585 560 798 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=102460 $D=1
M708 588 551 586 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=97830 $D=1
M709 589 552 587 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=102460 $D=1
M710 586 559 588 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=97830 $D=1
M711 587 560 589 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=102460 $D=1
M712 5 584 586 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=97830 $D=1
M713 6 585 587 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=102460 $D=1
M714 590 121 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=97830 $D=1
M715 591 121 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=102460 $D=1
M716 592 590 578 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=97830 $D=1
M717 593 591 579 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=102460 $D=1
M718 582 121 592 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=97830 $D=1
M719 583 121 593 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=102460 $D=1
M720 594 590 580 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=97830 $D=1
M721 595 591 581 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=102460 $D=1
M722 588 121 594 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=97830 $D=1
M723 589 121 595 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=102460 $D=1
M724 596 122 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=97830 $D=1
M725 597 122 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=102460 $D=1
M726 598 596 594 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=97830 $D=1
M727 599 597 595 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=102460 $D=1
M728 592 122 598 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=97830 $D=1
M729 593 122 599 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=102460 $D=1
M730 12 598 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=97830 $D=1
M731 13 599 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=102460 $D=1
M732 600 123 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=97830 $D=1
M733 601 123 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=102460 $D=1
M734 602 600 124 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=97830 $D=1
M735 603 601 125 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=102460 $D=1
M736 126 123 602 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=97830 $D=1
M737 127 123 603 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=102460 $D=1
M738 604 123 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=97830 $D=1
M739 605 123 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=102460 $D=1
M740 611 604 128 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=97830 $D=1
M741 612 605 130 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=102460 $D=1
M742 131 123 611 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=97830 $D=1
M743 129 123 612 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=102460 $D=1
M744 613 123 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=97830 $D=1
M745 614 123 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=102460 $D=1
M746 134 613 132 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=97830 $D=1
M747 134 614 133 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=102460 $D=1
M748 135 123 134 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=97830 $D=1
M749 136 123 134 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=102460 $D=1
M750 615 123 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=97830 $D=1
M751 616 123 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=102460 $D=1
M752 617 615 137 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=97830 $D=1
M753 618 616 138 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=102460 $D=1
M754 139 123 617 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=97830 $D=1
M755 140 123 618 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=102460 $D=1
M756 619 123 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=97830 $D=1
M757 620 123 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=102460 $D=1
M758 621 619 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=97830 $D=1
M759 622 620 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=102460 $D=1
M760 141 123 621 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=97830 $D=1
M761 142 123 622 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=102460 $D=1
M762 5 551 777 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=97830 $D=1
M763 6 552 778 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=102460 $D=1
M764 127 777 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=97830 $D=1
M765 124 778 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=102460 $D=1
M766 623 143 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=97830 $D=1
M767 624 143 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=102460 $D=1
M768 144 623 127 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=97830 $D=1
M769 145 624 124 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=102460 $D=1
M770 602 143 144 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=97830 $D=1
M771 603 143 145 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=102460 $D=1
M772 625 146 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=97830 $D=1
M773 626 146 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=102460 $D=1
M774 147 625 144 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=97830 $D=1
M775 148 626 145 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=102460 $D=1
M776 611 146 147 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=97830 $D=1
M777 612 146 148 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=102460 $D=1
M778 627 149 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=97830 $D=1
M779 628 149 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=102460 $D=1
M780 134 627 147 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=97830 $D=1
M781 150 628 148 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=102460 $D=1
M782 134 149 134 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=97830 $D=1
M783 134 149 150 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=102460 $D=1
M784 629 151 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=97830 $D=1
M785 630 151 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=102460 $D=1
M786 152 629 134 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=97830 $D=1
M787 153 630 150 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=102460 $D=1
M788 617 151 152 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=97830 $D=1
M789 618 151 153 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=102460 $D=1
M790 631 154 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=97830 $D=1
M791 632 154 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=102460 $D=1
M792 201 631 152 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=97830 $D=1
M793 202 632 153 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=102460 $D=1
M794 621 154 201 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=97830 $D=1
M795 622 154 202 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=102460 $D=1
M796 633 155 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=97830 $D=1
M797 634 155 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=102460 $D=1
M798 635 633 112 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=97830 $D=1
M799 636 634 113 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=102460 $D=1
M800 10 155 635 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=97830 $D=1
M801 11 155 636 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=102460 $D=1
M802 799 541 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=97830 $D=1
M803 800 542 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=102460 $D=1
M804 637 635 799 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=97830 $D=1
M805 638 636 800 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=102460 $D=1
M806 641 541 639 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=97830 $D=1
M807 642 542 640 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=102460 $D=1
M808 639 635 641 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=97830 $D=1
M809 640 636 642 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=102460 $D=1
M810 5 637 639 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=97830 $D=1
M811 6 638 640 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=102460 $D=1
M812 801 643 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=97830 $D=1
M813 802 644 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=102460 $D=1
M814 779 641 801 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=97830 $D=1
M815 780 642 802 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=102460 $D=1
M816 644 779 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=97830 $D=1
M817 156 780 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=102460 $D=1
M818 645 541 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=97830 $D=1
M819 646 542 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=102460 $D=1
M820 5 647 645 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=97830 $D=1
M821 6 648 646 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=102460 $D=1
M822 647 635 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=97830 $D=1
M823 648 636 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=102460 $D=1
M824 803 645 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=97830 $D=1
M825 804 646 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=102460 $D=1
M826 649 643 803 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=97830 $D=1
M827 650 644 804 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=102460 $D=1
M828 652 157 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=97830 $D=1
M829 653 651 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=102460 $D=1
M830 805 649 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=97830 $D=1
M831 806 650 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=102460 $D=1
M832 651 652 805 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=97830 $D=1
M833 158 653 806 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=102460 $D=1
M834 655 654 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=97830 $D=1
M835 656 159 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=102460 $D=1
M836 5 659 657 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=97830 $D=1
M837 6 660 658 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=102460 $D=1
M838 661 115 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=97830 $D=1
M839 662 116 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=102460 $D=1
M840 659 661 654 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=97830 $D=1
M841 660 662 159 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=102460 $D=1
M842 655 115 659 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=97830 $D=1
M843 656 116 660 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=102460 $D=1
M844 663 657 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=97830 $D=1
M845 664 658 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=102460 $D=1
M846 160 663 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=97830 $D=1
M847 654 664 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=102460 $D=1
M848 115 657 160 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=97830 $D=1
M849 116 658 654 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=102460 $D=1
M850 665 160 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=97830 $D=1
M851 666 654 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=102460 $D=1
M852 667 657 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=97830 $D=1
M853 668 658 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=102460 $D=1
M854 203 667 665 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=97830 $D=1
M855 204 668 666 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=102460 $D=1
M856 5 657 203 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=97830 $D=1
M857 6 658 204 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=102460 $D=1
M858 669 161 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=97830 $D=1
M859 670 161 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=102460 $D=1
M860 671 669 203 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=97830 $D=1
M861 672 670 204 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=102460 $D=1
M862 12 161 671 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=97830 $D=1
M863 13 161 672 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=102460 $D=1
M864 673 162 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=97830 $D=1
M865 674 162 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=102460 $D=1
M866 162 673 671 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=97830 $D=1
M867 162 674 672 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=102460 $D=1
M868 5 162 162 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=97830 $D=1
M869 6 162 162 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=102460 $D=1
M870 675 111 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=97830 $D=1
M871 676 111 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=102460 $D=1
M872 5 675 677 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=97830 $D=1
M873 6 676 678 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=102460 $D=1
M874 679 111 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=97830 $D=1
M875 680 111 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=102460 $D=1
M876 681 675 162 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=97830 $D=1
M877 682 676 162 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=102460 $D=1
M878 5 681 781 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=97830 $D=1
M879 6 682 782 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=102460 $D=1
M880 683 781 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=97830 $D=1
M881 684 782 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=102460 $D=1
M882 681 677 683 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=97830 $D=1
M883 682 678 684 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=102460 $D=1
M884 685 111 683 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=97830 $D=1
M885 686 111 684 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=102460 $D=1
M886 5 689 687 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=97830 $D=1
M887 6 690 688 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=102460 $D=1
M888 689 111 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=97830 $D=1
M889 690 111 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=102460 $D=1
M890 783 685 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=97830 $D=1
M891 784 686 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=102460 $D=1
M892 691 687 783 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=97830 $D=1
M893 692 688 784 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=102460 $D=1
M894 5 691 115 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=97830 $D=1
M895 6 692 116 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=102460 $D=1
M896 785 115 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=97830 $D=1
M897 786 116 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=102460 $D=1
M898 691 689 785 5 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=97830 $D=1
M899 692 690 786 6 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=102460 $D=1
M900 177 1 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=99080 $D=0
M901 178 1 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=103710 $D=0
M902 179 1 2 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=99080 $D=0
M903 180 1 3 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=103710 $D=0
M904 5 177 179 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=99080 $D=0
M905 6 178 180 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=103710 $D=0
M906 181 1 4 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=99080 $D=0
M907 182 1 4 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=103710 $D=0
M908 2 177 181 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=99080 $D=0
M909 3 178 182 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=103710 $D=0
M910 183 1 5 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=99080 $D=0
M911 184 1 6 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=103710 $D=0
M912 2 177 183 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=99080 $D=0
M913 3 178 184 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=103710 $D=0
M914 187 7 183 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=99080 $D=0
M915 188 7 184 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=103710 $D=0
M916 185 7 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=99080 $D=0
M917 186 7 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=103710 $D=0
M918 189 7 181 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=99080 $D=0
M919 190 7 182 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=103710 $D=0
M920 179 185 189 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=99080 $D=0
M921 180 186 190 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=103710 $D=0
M922 191 8 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=99080 $D=0
M923 192 8 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=103710 $D=0
M924 193 8 189 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=99080 $D=0
M925 194 8 190 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=103710 $D=0
M926 187 191 193 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=99080 $D=0
M927 188 192 194 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=103710 $D=0
M928 195 9 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=99080 $D=0
M929 196 9 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=103710 $D=0
M930 197 9 5 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=99080 $D=0
M931 198 9 6 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=103710 $D=0
M932 10 195 197 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=99080 $D=0
M933 11 196 198 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=103710 $D=0
M934 199 9 12 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=99080 $D=0
M935 200 9 13 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=103710 $D=0
M936 201 195 199 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=99080 $D=0
M937 202 196 200 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=103710 $D=0
M938 205 9 203 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=99080 $D=0
M939 206 9 204 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=103710 $D=0
M940 193 195 205 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=99080 $D=0
M941 194 196 206 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=103710 $D=0
M942 209 14 205 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=99080 $D=0
M943 210 14 206 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=103710 $D=0
M944 207 14 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=99080 $D=0
M945 208 14 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=103710 $D=0
M946 211 14 199 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=99080 $D=0
M947 212 14 200 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=103710 $D=0
M948 197 207 211 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=99080 $D=0
M949 198 208 212 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=103710 $D=0
M950 213 15 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=99080 $D=0
M951 214 15 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=103710 $D=0
M952 215 15 211 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=99080 $D=0
M953 216 15 212 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=103710 $D=0
M954 209 213 215 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=99080 $D=0
M955 210 214 216 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=103710 $D=0
M956 163 16 217 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=99080 $D=0
M957 164 16 218 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=103710 $D=0
M958 219 17 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=99080 $D=0
M959 220 17 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=103710 $D=0
M960 221 217 215 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=99080 $D=0
M961 222 218 216 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=103710 $D=0
M962 163 221 693 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=99080 $D=0
M963 164 222 694 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=103710 $D=0
M964 223 693 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=99080 $D=0
M965 224 694 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=103710 $D=0
M966 221 16 223 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=99080 $D=0
M967 222 16 224 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=103710 $D=0
M968 223 219 225 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=99080 $D=0
M969 224 220 226 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=103710 $D=0
M970 229 227 223 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=99080 $D=0
M971 230 228 224 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=103710 $D=0
M972 227 18 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=99080 $D=0
M973 228 18 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=103710 $D=0
M974 163 19 231 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=99080 $D=0
M975 164 19 232 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=103710 $D=0
M976 233 20 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=99080 $D=0
M977 234 20 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=103710 $D=0
M978 235 231 215 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=99080 $D=0
M979 236 232 216 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=103710 $D=0
M980 163 235 695 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=99080 $D=0
M981 164 236 696 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=103710 $D=0
M982 237 695 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=99080 $D=0
M983 238 696 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=103710 $D=0
M984 235 19 237 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=99080 $D=0
M985 236 19 238 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=103710 $D=0
M986 237 233 225 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=99080 $D=0
M987 238 234 226 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=103710 $D=0
M988 229 239 237 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=99080 $D=0
M989 230 240 238 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=103710 $D=0
M990 239 21 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=99080 $D=0
M991 240 21 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=103710 $D=0
M992 163 22 241 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=99080 $D=0
M993 164 22 242 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=103710 $D=0
M994 243 23 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=99080 $D=0
M995 244 23 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=103710 $D=0
M996 245 241 215 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=99080 $D=0
M997 246 242 216 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=103710 $D=0
M998 163 245 697 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=99080 $D=0
M999 164 246 698 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=103710 $D=0
M1000 247 697 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=99080 $D=0
M1001 248 698 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=103710 $D=0
M1002 245 22 247 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=99080 $D=0
M1003 246 22 248 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=103710 $D=0
M1004 247 243 225 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=99080 $D=0
M1005 248 244 226 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=103710 $D=0
M1006 229 249 247 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=99080 $D=0
M1007 230 250 248 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=103710 $D=0
M1008 249 24 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=99080 $D=0
M1009 250 24 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=103710 $D=0
M1010 163 25 251 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=99080 $D=0
M1011 164 25 252 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=103710 $D=0
M1012 253 26 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=99080 $D=0
M1013 254 26 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=103710 $D=0
M1014 255 251 215 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=99080 $D=0
M1015 256 252 216 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=103710 $D=0
M1016 163 255 699 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=99080 $D=0
M1017 164 256 700 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=103710 $D=0
M1018 257 699 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=99080 $D=0
M1019 258 700 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=103710 $D=0
M1020 255 25 257 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=99080 $D=0
M1021 256 25 258 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=103710 $D=0
M1022 257 253 225 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=99080 $D=0
M1023 258 254 226 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=103710 $D=0
M1024 229 259 257 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=99080 $D=0
M1025 230 260 258 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=103710 $D=0
M1026 259 27 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=99080 $D=0
M1027 260 27 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=103710 $D=0
M1028 163 28 261 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=99080 $D=0
M1029 164 28 262 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=103710 $D=0
M1030 263 29 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=99080 $D=0
M1031 264 29 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=103710 $D=0
M1032 265 261 215 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=99080 $D=0
M1033 266 262 216 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=103710 $D=0
M1034 163 265 701 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=99080 $D=0
M1035 164 266 702 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=103710 $D=0
M1036 267 701 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=99080 $D=0
M1037 268 702 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=103710 $D=0
M1038 265 28 267 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=99080 $D=0
M1039 266 28 268 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=103710 $D=0
M1040 267 263 225 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=99080 $D=0
M1041 268 264 226 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=103710 $D=0
M1042 229 269 267 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=99080 $D=0
M1043 230 270 268 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=103710 $D=0
M1044 269 30 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=99080 $D=0
M1045 270 30 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=103710 $D=0
M1046 163 31 271 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=99080 $D=0
M1047 164 31 272 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=103710 $D=0
M1048 273 32 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=99080 $D=0
M1049 274 32 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=103710 $D=0
M1050 275 271 215 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=99080 $D=0
M1051 276 272 216 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=103710 $D=0
M1052 163 275 703 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=99080 $D=0
M1053 164 276 704 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=103710 $D=0
M1054 277 703 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=99080 $D=0
M1055 278 704 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=103710 $D=0
M1056 275 31 277 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=99080 $D=0
M1057 276 31 278 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=103710 $D=0
M1058 277 273 225 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=99080 $D=0
M1059 278 274 226 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=103710 $D=0
M1060 229 279 277 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=99080 $D=0
M1061 230 280 278 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=103710 $D=0
M1062 279 33 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=99080 $D=0
M1063 280 33 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=103710 $D=0
M1064 163 34 281 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=99080 $D=0
M1065 164 34 282 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=103710 $D=0
M1066 283 35 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=99080 $D=0
M1067 284 35 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=103710 $D=0
M1068 285 281 215 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=99080 $D=0
M1069 286 282 216 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=103710 $D=0
M1070 163 285 705 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=99080 $D=0
M1071 164 286 706 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=103710 $D=0
M1072 287 705 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=99080 $D=0
M1073 288 706 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=103710 $D=0
M1074 285 34 287 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=99080 $D=0
M1075 286 34 288 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=103710 $D=0
M1076 287 283 225 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=99080 $D=0
M1077 288 284 226 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=103710 $D=0
M1078 229 289 287 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=99080 $D=0
M1079 230 290 288 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=103710 $D=0
M1080 289 36 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=99080 $D=0
M1081 290 36 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=103710 $D=0
M1082 163 37 291 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=99080 $D=0
M1083 164 37 292 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=103710 $D=0
M1084 293 38 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=99080 $D=0
M1085 294 38 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=103710 $D=0
M1086 295 291 215 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=99080 $D=0
M1087 296 292 216 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=103710 $D=0
M1088 163 295 707 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=99080 $D=0
M1089 164 296 708 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=103710 $D=0
M1090 297 707 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=99080 $D=0
M1091 298 708 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=103710 $D=0
M1092 295 37 297 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=99080 $D=0
M1093 296 37 298 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=103710 $D=0
M1094 297 293 225 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=99080 $D=0
M1095 298 294 226 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=103710 $D=0
M1096 229 299 297 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=99080 $D=0
M1097 230 300 298 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=103710 $D=0
M1098 299 39 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=99080 $D=0
M1099 300 39 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=103710 $D=0
M1100 163 40 301 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=99080 $D=0
M1101 164 40 302 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=103710 $D=0
M1102 303 41 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=99080 $D=0
M1103 304 41 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=103710 $D=0
M1104 305 301 215 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=99080 $D=0
M1105 306 302 216 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=103710 $D=0
M1106 163 305 709 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=99080 $D=0
M1107 164 306 710 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=103710 $D=0
M1108 307 709 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=99080 $D=0
M1109 308 710 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=103710 $D=0
M1110 305 40 307 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=99080 $D=0
M1111 306 40 308 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=103710 $D=0
M1112 307 303 225 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=99080 $D=0
M1113 308 304 226 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=103710 $D=0
M1114 229 309 307 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=99080 $D=0
M1115 230 310 308 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=103710 $D=0
M1116 309 42 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=99080 $D=0
M1117 310 42 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=103710 $D=0
M1118 163 43 311 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=99080 $D=0
M1119 164 43 312 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=103710 $D=0
M1120 313 44 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=99080 $D=0
M1121 314 44 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=103710 $D=0
M1122 315 311 215 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=99080 $D=0
M1123 316 312 216 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=103710 $D=0
M1124 163 315 711 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=99080 $D=0
M1125 164 316 712 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=103710 $D=0
M1126 317 711 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=99080 $D=0
M1127 318 712 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=103710 $D=0
M1128 315 43 317 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=99080 $D=0
M1129 316 43 318 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=103710 $D=0
M1130 317 313 225 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=99080 $D=0
M1131 318 314 226 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=103710 $D=0
M1132 229 319 317 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=99080 $D=0
M1133 230 320 318 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=103710 $D=0
M1134 319 45 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=99080 $D=0
M1135 320 45 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=103710 $D=0
M1136 163 46 321 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=99080 $D=0
M1137 164 46 322 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=103710 $D=0
M1138 323 47 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=99080 $D=0
M1139 324 47 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=103710 $D=0
M1140 325 321 215 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=99080 $D=0
M1141 326 322 216 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=103710 $D=0
M1142 163 325 713 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=99080 $D=0
M1143 164 326 714 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=103710 $D=0
M1144 327 713 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=99080 $D=0
M1145 328 714 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=103710 $D=0
M1146 325 46 327 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=99080 $D=0
M1147 326 46 328 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=103710 $D=0
M1148 327 323 225 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=99080 $D=0
M1149 328 324 226 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=103710 $D=0
M1150 229 329 327 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=99080 $D=0
M1151 230 330 328 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=103710 $D=0
M1152 329 48 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=99080 $D=0
M1153 330 48 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=103710 $D=0
M1154 163 49 331 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=99080 $D=0
M1155 164 49 332 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=103710 $D=0
M1156 333 50 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=99080 $D=0
M1157 334 50 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=103710 $D=0
M1158 335 331 215 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=99080 $D=0
M1159 336 332 216 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=103710 $D=0
M1160 163 335 715 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=99080 $D=0
M1161 164 336 716 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=103710 $D=0
M1162 337 715 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=99080 $D=0
M1163 338 716 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=103710 $D=0
M1164 335 49 337 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=99080 $D=0
M1165 336 49 338 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=103710 $D=0
M1166 337 333 225 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=99080 $D=0
M1167 338 334 226 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=103710 $D=0
M1168 229 339 337 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=99080 $D=0
M1169 230 340 338 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=103710 $D=0
M1170 339 51 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=99080 $D=0
M1171 340 51 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=103710 $D=0
M1172 163 52 341 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=99080 $D=0
M1173 164 52 342 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=103710 $D=0
M1174 343 53 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=99080 $D=0
M1175 344 53 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=103710 $D=0
M1176 345 341 215 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=99080 $D=0
M1177 346 342 216 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=103710 $D=0
M1178 163 345 717 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=99080 $D=0
M1179 164 346 718 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=103710 $D=0
M1180 347 717 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=99080 $D=0
M1181 348 718 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=103710 $D=0
M1182 345 52 347 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=99080 $D=0
M1183 346 52 348 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=103710 $D=0
M1184 347 343 225 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=99080 $D=0
M1185 348 344 226 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=103710 $D=0
M1186 229 349 347 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=99080 $D=0
M1187 230 350 348 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=103710 $D=0
M1188 349 54 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=99080 $D=0
M1189 350 54 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=103710 $D=0
M1190 163 55 351 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=99080 $D=0
M1191 164 55 352 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=103710 $D=0
M1192 353 56 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=99080 $D=0
M1193 354 56 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=103710 $D=0
M1194 355 351 215 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=99080 $D=0
M1195 356 352 216 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=103710 $D=0
M1196 163 355 719 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=99080 $D=0
M1197 164 356 720 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=103710 $D=0
M1198 357 719 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=99080 $D=0
M1199 358 720 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=103710 $D=0
M1200 355 55 357 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=99080 $D=0
M1201 356 55 358 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=103710 $D=0
M1202 357 353 225 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=99080 $D=0
M1203 358 354 226 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=103710 $D=0
M1204 229 359 357 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=99080 $D=0
M1205 230 360 358 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=103710 $D=0
M1206 359 57 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=99080 $D=0
M1207 360 57 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=103710 $D=0
M1208 163 58 361 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=99080 $D=0
M1209 164 58 362 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=103710 $D=0
M1210 363 59 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=99080 $D=0
M1211 364 59 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=103710 $D=0
M1212 365 361 215 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=99080 $D=0
M1213 366 362 216 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=103710 $D=0
M1214 163 365 721 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=99080 $D=0
M1215 164 366 722 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=103710 $D=0
M1216 367 721 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=99080 $D=0
M1217 368 722 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=103710 $D=0
M1218 365 58 367 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=99080 $D=0
M1219 366 58 368 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=103710 $D=0
M1220 367 363 225 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=99080 $D=0
M1221 368 364 226 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=103710 $D=0
M1222 229 369 367 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=99080 $D=0
M1223 230 370 368 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=103710 $D=0
M1224 369 60 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=99080 $D=0
M1225 370 60 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=103710 $D=0
M1226 163 61 371 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=99080 $D=0
M1227 164 61 372 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=103710 $D=0
M1228 373 62 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=99080 $D=0
M1229 374 62 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=103710 $D=0
M1230 375 371 215 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=99080 $D=0
M1231 376 372 216 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=103710 $D=0
M1232 163 375 723 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=99080 $D=0
M1233 164 376 724 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=103710 $D=0
M1234 377 723 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=99080 $D=0
M1235 378 724 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=103710 $D=0
M1236 375 61 377 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=99080 $D=0
M1237 376 61 378 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=103710 $D=0
M1238 377 373 225 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=99080 $D=0
M1239 378 374 226 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=103710 $D=0
M1240 229 379 377 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=99080 $D=0
M1241 230 380 378 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=103710 $D=0
M1242 379 63 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=99080 $D=0
M1243 380 63 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=103710 $D=0
M1244 163 64 381 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=99080 $D=0
M1245 164 64 382 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=103710 $D=0
M1246 383 65 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=99080 $D=0
M1247 384 65 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=103710 $D=0
M1248 385 381 215 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=99080 $D=0
M1249 386 382 216 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=103710 $D=0
M1250 163 385 725 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=99080 $D=0
M1251 164 386 726 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=103710 $D=0
M1252 387 725 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=99080 $D=0
M1253 388 726 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=103710 $D=0
M1254 385 64 387 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=99080 $D=0
M1255 386 64 388 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=103710 $D=0
M1256 387 383 225 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=99080 $D=0
M1257 388 384 226 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=103710 $D=0
M1258 229 389 387 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=99080 $D=0
M1259 230 390 388 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=103710 $D=0
M1260 389 66 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=99080 $D=0
M1261 390 66 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=103710 $D=0
M1262 163 67 391 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=99080 $D=0
M1263 164 67 392 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=103710 $D=0
M1264 393 68 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=99080 $D=0
M1265 394 68 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=103710 $D=0
M1266 395 391 215 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=99080 $D=0
M1267 396 392 216 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=103710 $D=0
M1268 163 395 727 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=99080 $D=0
M1269 164 396 728 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=103710 $D=0
M1270 397 727 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=99080 $D=0
M1271 398 728 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=103710 $D=0
M1272 395 67 397 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=99080 $D=0
M1273 396 67 398 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=103710 $D=0
M1274 397 393 225 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=99080 $D=0
M1275 398 394 226 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=103710 $D=0
M1276 229 399 397 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=99080 $D=0
M1277 230 400 398 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=103710 $D=0
M1278 399 69 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=99080 $D=0
M1279 400 69 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=103710 $D=0
M1280 163 70 401 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=99080 $D=0
M1281 164 70 402 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=103710 $D=0
M1282 403 71 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=99080 $D=0
M1283 404 71 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=103710 $D=0
M1284 405 401 215 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=99080 $D=0
M1285 406 402 216 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=103710 $D=0
M1286 163 405 729 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=99080 $D=0
M1287 164 406 730 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=103710 $D=0
M1288 407 729 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=99080 $D=0
M1289 408 730 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=103710 $D=0
M1290 405 70 407 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=99080 $D=0
M1291 406 70 408 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=103710 $D=0
M1292 407 403 225 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=99080 $D=0
M1293 408 404 226 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=103710 $D=0
M1294 229 409 407 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=99080 $D=0
M1295 230 410 408 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=103710 $D=0
M1296 409 72 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=99080 $D=0
M1297 410 72 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=103710 $D=0
M1298 163 73 411 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=99080 $D=0
M1299 164 73 412 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=103710 $D=0
M1300 413 74 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=99080 $D=0
M1301 414 74 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=103710 $D=0
M1302 415 411 215 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=99080 $D=0
M1303 416 412 216 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=103710 $D=0
M1304 163 415 731 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=99080 $D=0
M1305 164 416 732 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=103710 $D=0
M1306 417 731 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=99080 $D=0
M1307 418 732 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=103710 $D=0
M1308 415 73 417 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=99080 $D=0
M1309 416 73 418 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=103710 $D=0
M1310 417 413 225 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=99080 $D=0
M1311 418 414 226 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=103710 $D=0
M1312 229 419 417 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=99080 $D=0
M1313 230 420 418 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=103710 $D=0
M1314 419 75 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=99080 $D=0
M1315 420 75 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=103710 $D=0
M1316 163 76 421 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=99080 $D=0
M1317 164 76 422 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=103710 $D=0
M1318 423 77 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=99080 $D=0
M1319 424 77 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=103710 $D=0
M1320 425 421 215 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=99080 $D=0
M1321 426 422 216 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=103710 $D=0
M1322 163 425 733 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=99080 $D=0
M1323 164 426 734 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=103710 $D=0
M1324 427 733 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=99080 $D=0
M1325 428 734 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=103710 $D=0
M1326 425 76 427 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=99080 $D=0
M1327 426 76 428 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=103710 $D=0
M1328 427 423 225 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=99080 $D=0
M1329 428 424 226 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=103710 $D=0
M1330 229 429 427 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=99080 $D=0
M1331 230 430 428 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=103710 $D=0
M1332 429 78 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=99080 $D=0
M1333 430 78 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=103710 $D=0
M1334 163 79 431 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=99080 $D=0
M1335 164 79 432 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=103710 $D=0
M1336 433 80 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=99080 $D=0
M1337 434 80 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=103710 $D=0
M1338 435 431 215 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=99080 $D=0
M1339 436 432 216 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=103710 $D=0
M1340 163 435 735 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=99080 $D=0
M1341 164 436 736 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=103710 $D=0
M1342 437 735 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=99080 $D=0
M1343 438 736 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=103710 $D=0
M1344 435 79 437 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=99080 $D=0
M1345 436 79 438 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=103710 $D=0
M1346 437 433 225 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=99080 $D=0
M1347 438 434 226 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=103710 $D=0
M1348 229 439 437 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=99080 $D=0
M1349 230 440 438 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=103710 $D=0
M1350 439 81 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=99080 $D=0
M1351 440 81 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=103710 $D=0
M1352 163 82 441 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=99080 $D=0
M1353 164 82 442 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=103710 $D=0
M1354 443 83 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=99080 $D=0
M1355 444 83 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=103710 $D=0
M1356 445 441 215 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=99080 $D=0
M1357 446 442 216 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=103710 $D=0
M1358 163 445 737 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=99080 $D=0
M1359 164 446 738 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=103710 $D=0
M1360 447 737 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=99080 $D=0
M1361 448 738 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=103710 $D=0
M1362 445 82 447 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=99080 $D=0
M1363 446 82 448 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=103710 $D=0
M1364 447 443 225 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=99080 $D=0
M1365 448 444 226 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=103710 $D=0
M1366 229 449 447 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=99080 $D=0
M1367 230 450 448 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=103710 $D=0
M1368 449 84 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=99080 $D=0
M1369 450 84 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=103710 $D=0
M1370 163 85 451 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=99080 $D=0
M1371 164 85 452 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=103710 $D=0
M1372 453 86 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=99080 $D=0
M1373 454 86 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=103710 $D=0
M1374 455 451 215 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=99080 $D=0
M1375 456 452 216 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=103710 $D=0
M1376 163 455 739 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=99080 $D=0
M1377 164 456 740 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=103710 $D=0
M1378 457 739 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=99080 $D=0
M1379 458 740 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=103710 $D=0
M1380 455 85 457 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=99080 $D=0
M1381 456 85 458 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=103710 $D=0
M1382 457 453 225 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=99080 $D=0
M1383 458 454 226 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=103710 $D=0
M1384 229 459 457 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=99080 $D=0
M1385 230 460 458 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=103710 $D=0
M1386 459 87 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=99080 $D=0
M1387 460 87 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=103710 $D=0
M1388 163 88 461 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=99080 $D=0
M1389 164 88 462 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=103710 $D=0
M1390 463 89 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=99080 $D=0
M1391 464 89 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=103710 $D=0
M1392 465 461 215 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=99080 $D=0
M1393 466 462 216 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=103710 $D=0
M1394 163 465 741 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=99080 $D=0
M1395 164 466 742 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=103710 $D=0
M1396 467 741 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=99080 $D=0
M1397 468 742 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=103710 $D=0
M1398 465 88 467 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=99080 $D=0
M1399 466 88 468 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=103710 $D=0
M1400 467 463 225 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=99080 $D=0
M1401 468 464 226 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=103710 $D=0
M1402 229 469 467 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=99080 $D=0
M1403 230 470 468 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=103710 $D=0
M1404 469 90 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=99080 $D=0
M1405 470 90 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=103710 $D=0
M1406 163 91 471 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=99080 $D=0
M1407 164 91 472 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=103710 $D=0
M1408 473 92 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=99080 $D=0
M1409 474 92 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=103710 $D=0
M1410 475 471 215 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=99080 $D=0
M1411 476 472 216 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=103710 $D=0
M1412 163 475 743 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=99080 $D=0
M1413 164 476 744 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=103710 $D=0
M1414 477 743 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=99080 $D=0
M1415 478 744 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=103710 $D=0
M1416 475 91 477 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=99080 $D=0
M1417 476 91 478 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=103710 $D=0
M1418 477 473 225 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=99080 $D=0
M1419 478 474 226 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=103710 $D=0
M1420 229 479 477 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=99080 $D=0
M1421 230 480 478 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=103710 $D=0
M1422 479 93 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=99080 $D=0
M1423 480 93 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=103710 $D=0
M1424 163 94 481 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=99080 $D=0
M1425 164 94 482 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=103710 $D=0
M1426 483 95 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=99080 $D=0
M1427 484 95 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=103710 $D=0
M1428 485 481 215 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=99080 $D=0
M1429 486 482 216 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=103710 $D=0
M1430 163 485 745 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=99080 $D=0
M1431 164 486 746 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=103710 $D=0
M1432 487 745 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=99080 $D=0
M1433 488 746 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=103710 $D=0
M1434 485 94 487 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=99080 $D=0
M1435 486 94 488 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=103710 $D=0
M1436 487 483 225 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=99080 $D=0
M1437 488 484 226 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=103710 $D=0
M1438 229 489 487 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=99080 $D=0
M1439 230 490 488 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=103710 $D=0
M1440 489 96 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=99080 $D=0
M1441 490 96 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=103710 $D=0
M1442 163 97 491 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=99080 $D=0
M1443 164 97 492 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=103710 $D=0
M1444 493 98 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=99080 $D=0
M1445 494 98 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=103710 $D=0
M1446 495 491 215 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=99080 $D=0
M1447 496 492 216 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=103710 $D=0
M1448 163 495 747 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=99080 $D=0
M1449 164 496 748 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=103710 $D=0
M1450 497 747 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=99080 $D=0
M1451 498 748 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=103710 $D=0
M1452 495 97 497 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=99080 $D=0
M1453 496 97 498 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=103710 $D=0
M1454 497 493 225 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=99080 $D=0
M1455 498 494 226 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=103710 $D=0
M1456 229 499 497 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=99080 $D=0
M1457 230 500 498 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=103710 $D=0
M1458 499 99 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=99080 $D=0
M1459 500 99 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=103710 $D=0
M1460 163 100 501 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=99080 $D=0
M1461 164 100 502 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=103710 $D=0
M1462 503 101 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=99080 $D=0
M1463 504 101 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=103710 $D=0
M1464 505 501 215 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=99080 $D=0
M1465 506 502 216 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=103710 $D=0
M1466 163 505 749 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=99080 $D=0
M1467 164 506 750 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=103710 $D=0
M1468 507 749 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=99080 $D=0
M1469 508 750 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=103710 $D=0
M1470 505 100 507 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=99080 $D=0
M1471 506 100 508 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=103710 $D=0
M1472 507 503 225 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=99080 $D=0
M1473 508 504 226 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=103710 $D=0
M1474 229 509 507 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=99080 $D=0
M1475 230 510 508 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=103710 $D=0
M1476 509 102 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=99080 $D=0
M1477 510 102 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=103710 $D=0
M1478 163 103 511 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=99080 $D=0
M1479 164 103 512 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=103710 $D=0
M1480 513 104 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=99080 $D=0
M1481 514 104 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=103710 $D=0
M1482 515 511 215 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=99080 $D=0
M1483 516 512 216 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=103710 $D=0
M1484 163 515 751 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=99080 $D=0
M1485 164 516 752 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=103710 $D=0
M1486 517 751 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=99080 $D=0
M1487 518 752 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=103710 $D=0
M1488 515 103 517 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=99080 $D=0
M1489 516 103 518 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=103710 $D=0
M1490 517 513 225 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=99080 $D=0
M1491 518 514 226 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=103710 $D=0
M1492 229 519 517 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=99080 $D=0
M1493 230 520 518 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=103710 $D=0
M1494 519 105 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=99080 $D=0
M1495 520 105 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=103710 $D=0
M1496 163 106 521 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=99080 $D=0
M1497 164 106 522 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=103710 $D=0
M1498 523 107 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=99080 $D=0
M1499 524 107 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=103710 $D=0
M1500 525 521 215 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=99080 $D=0
M1501 526 522 216 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=103710 $D=0
M1502 163 525 753 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=99080 $D=0
M1503 164 526 754 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=103710 $D=0
M1504 527 753 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=99080 $D=0
M1505 528 754 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=103710 $D=0
M1506 525 106 527 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=99080 $D=0
M1507 526 106 528 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=103710 $D=0
M1508 527 523 225 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=99080 $D=0
M1509 528 524 226 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=103710 $D=0
M1510 229 529 527 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=99080 $D=0
M1511 230 530 528 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=103710 $D=0
M1512 529 108 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=99080 $D=0
M1513 530 108 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=103710 $D=0
M1514 163 109 531 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=99080 $D=0
M1515 164 109 532 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=103710 $D=0
M1516 533 110 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=99080 $D=0
M1517 534 110 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=103710 $D=0
M1518 5 533 225 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=99080 $D=0
M1519 6 534 226 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=103710 $D=0
M1520 229 531 5 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=99080 $D=0
M1521 230 532 6 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=103710 $D=0
M1522 163 537 535 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=99080 $D=0
M1523 164 538 536 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=103710 $D=0
M1524 537 111 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=99080 $D=0
M1525 538 111 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=103710 $D=0
M1526 755 225 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=99080 $D=0
M1527 756 226 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=103710 $D=0
M1528 539 537 755 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=99080 $D=0
M1529 540 538 756 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=103710 $D=0
M1530 163 539 541 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=99080 $D=0
M1531 164 540 542 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=103710 $D=0
M1532 757 541 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=99080 $D=0
M1533 758 542 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=103710 $D=0
M1534 539 535 757 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=99080 $D=0
M1535 540 536 758 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=103710 $D=0
M1536 163 545 543 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=99080 $D=0
M1537 164 546 544 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=103710 $D=0
M1538 545 111 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=99080 $D=0
M1539 546 111 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=103710 $D=0
M1540 759 229 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=99080 $D=0
M1541 760 230 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=103710 $D=0
M1542 547 545 759 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=99080 $D=0
M1543 548 546 760 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=103710 $D=0
M1544 163 547 112 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=99080 $D=0
M1545 164 548 113 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=103710 $D=0
M1546 761 112 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=99080 $D=0
M1547 762 113 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=103710 $D=0
M1548 547 543 761 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=99080 $D=0
M1549 548 544 762 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=103710 $D=0
M1550 549 114 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=99080 $D=0
M1551 550 114 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=103710 $D=0
M1552 551 114 541 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=99080 $D=0
M1553 552 114 542 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=103710 $D=0
M1554 115 549 551 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=99080 $D=0
M1555 116 550 552 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=103710 $D=0
M1556 553 117 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=99080 $D=0
M1557 554 117 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=103710 $D=0
M1558 555 117 112 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=99080 $D=0
M1559 556 117 113 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=103710 $D=0
M1560 763 553 555 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=99080 $D=0
M1561 764 554 556 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=103710 $D=0
M1562 163 112 763 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=99080 $D=0
M1563 164 113 764 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=103710 $D=0
M1564 557 118 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=99080 $D=0
M1565 558 118 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=103710 $D=0
M1566 559 118 555 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=99080 $D=0
M1567 560 118 556 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=103710 $D=0
M1568 10 557 559 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=99080 $D=0
M1569 11 558 560 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=103710 $D=0
M1570 562 561 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=99080 $D=0
M1571 563 119 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=103710 $D=0
M1572 163 566 564 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=99080 $D=0
M1573 164 567 565 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=103710 $D=0
M1574 568 551 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=99080 $D=0
M1575 569 552 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=103710 $D=0
M1576 566 551 561 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=99080 $D=0
M1577 567 552 119 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=103710 $D=0
M1578 562 568 566 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=99080 $D=0
M1579 563 569 567 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=103710 $D=0
M1580 570 564 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=99080 $D=0
M1581 571 565 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=103710 $D=0
M1582 120 564 559 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=99080 $D=0
M1583 561 565 560 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=103710 $D=0
M1584 551 570 120 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=99080 $D=0
M1585 552 571 561 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=103710 $D=0
M1586 572 120 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=99080 $D=0
M1587 573 561 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=103710 $D=0
M1588 574 564 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=99080 $D=0
M1589 575 565 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=103710 $D=0
M1590 576 564 572 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=99080 $D=0
M1591 577 565 573 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=103710 $D=0
M1592 559 574 576 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=99080 $D=0
M1593 560 575 577 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=103710 $D=0
M1594 787 551 163 163 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=98720 $D=0
M1595 788 552 164 164 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=103350 $D=0
M1596 578 559 787 163 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=98720 $D=0
M1597 579 560 788 164 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=103350 $D=0
M1598 580 576 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=99080 $D=0
M1599 581 577 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=103710 $D=0
M1600 582 551 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=99080 $D=0
M1601 583 552 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=103710 $D=0
M1602 163 559 582 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=99080 $D=0
M1603 164 560 583 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=103710 $D=0
M1604 584 551 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=99080 $D=0
M1605 585 552 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=103710 $D=0
M1606 163 559 584 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=99080 $D=0
M1607 164 560 585 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=103710 $D=0
M1608 789 551 163 163 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=98900 $D=0
M1609 790 552 164 164 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=103530 $D=0
M1610 588 559 789 163 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=98900 $D=0
M1611 589 560 790 164 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=103530 $D=0
M1612 163 584 588 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=99080 $D=0
M1613 164 585 589 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=103710 $D=0
M1614 590 121 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=99080 $D=0
M1615 591 121 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=103710 $D=0
M1616 592 121 578 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=99080 $D=0
M1617 593 121 579 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=103710 $D=0
M1618 582 590 592 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=99080 $D=0
M1619 583 591 593 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=103710 $D=0
M1620 594 121 580 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=99080 $D=0
M1621 595 121 581 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=103710 $D=0
M1622 588 590 594 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=99080 $D=0
M1623 589 591 595 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=103710 $D=0
M1624 596 122 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=99080 $D=0
M1625 597 122 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=103710 $D=0
M1626 598 122 594 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=99080 $D=0
M1627 599 122 595 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=103710 $D=0
M1628 592 596 598 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=99080 $D=0
M1629 593 597 599 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=103710 $D=0
M1630 12 598 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=99080 $D=0
M1631 13 599 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=103710 $D=0
M1632 600 123 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=99080 $D=0
M1633 601 123 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=103710 $D=0
M1634 602 123 124 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=99080 $D=0
M1635 603 123 125 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=103710 $D=0
M1636 126 600 602 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=99080 $D=0
M1637 127 601 603 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=103710 $D=0
M1638 604 123 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=99080 $D=0
M1639 605 123 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=103710 $D=0
M1640 611 123 128 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=99080 $D=0
M1641 612 123 130 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=103710 $D=0
M1642 131 604 611 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=99080 $D=0
M1643 129 605 612 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=103710 $D=0
M1644 613 123 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=99080 $D=0
M1645 614 123 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=103710 $D=0
M1646 134 123 132 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=99080 $D=0
M1647 134 123 133 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=103710 $D=0
M1648 135 613 134 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=99080 $D=0
M1649 136 614 134 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=103710 $D=0
M1650 615 123 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=99080 $D=0
M1651 616 123 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=103710 $D=0
M1652 617 123 137 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=99080 $D=0
M1653 618 123 138 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=103710 $D=0
M1654 139 615 617 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=99080 $D=0
M1655 140 616 618 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=103710 $D=0
M1656 619 123 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=99080 $D=0
M1657 620 123 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=103710 $D=0
M1658 621 123 5 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=99080 $D=0
M1659 622 123 6 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=103710 $D=0
M1660 141 619 621 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=99080 $D=0
M1661 142 620 622 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=103710 $D=0
M1662 163 551 777 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=99080 $D=0
M1663 164 552 778 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=103710 $D=0
M1664 127 777 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=99080 $D=0
M1665 124 778 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=103710 $D=0
M1666 623 143 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=99080 $D=0
M1667 624 143 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=103710 $D=0
M1668 144 143 127 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=99080 $D=0
M1669 145 143 124 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=103710 $D=0
M1670 602 623 144 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=99080 $D=0
M1671 603 624 145 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=103710 $D=0
M1672 625 146 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=99080 $D=0
M1673 626 146 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=103710 $D=0
M1674 147 146 144 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=99080 $D=0
M1675 148 146 145 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=103710 $D=0
M1676 611 625 147 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=99080 $D=0
M1677 612 626 148 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=103710 $D=0
M1678 627 149 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=99080 $D=0
M1679 628 149 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=103710 $D=0
M1680 134 149 147 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=99080 $D=0
M1681 150 149 148 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=103710 $D=0
M1682 134 627 134 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=99080 $D=0
M1683 134 628 150 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=103710 $D=0
M1684 629 151 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=99080 $D=0
M1685 630 151 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=103710 $D=0
M1686 152 151 134 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=99080 $D=0
M1687 153 151 150 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=103710 $D=0
M1688 617 629 152 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=99080 $D=0
M1689 618 630 153 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=103710 $D=0
M1690 631 154 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=99080 $D=0
M1691 632 154 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=103710 $D=0
M1692 201 154 152 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=99080 $D=0
M1693 202 154 153 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=103710 $D=0
M1694 621 631 201 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=99080 $D=0
M1695 622 632 202 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=103710 $D=0
M1696 633 155 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=99080 $D=0
M1697 634 155 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=103710 $D=0
M1698 635 155 112 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=99080 $D=0
M1699 636 155 113 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=103710 $D=0
M1700 10 633 635 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=99080 $D=0
M1701 11 634 636 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=103710 $D=0
M1702 637 541 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=99080 $D=0
M1703 638 542 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=103710 $D=0
M1704 163 635 637 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=99080 $D=0
M1705 164 636 638 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=103710 $D=0
M1706 791 541 163 163 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=98900 $D=0
M1707 792 542 164 164 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=103530 $D=0
M1708 641 635 791 163 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=98900 $D=0
M1709 642 636 792 164 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=103530 $D=0
M1710 163 637 641 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=99080 $D=0
M1711 164 638 642 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=103710 $D=0
M1712 779 643 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=99080 $D=0
M1713 780 644 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=103710 $D=0
M1714 163 641 779 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=99080 $D=0
M1715 164 642 780 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=103710 $D=0
M1716 644 779 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=99080 $D=0
M1717 156 780 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=103710 $D=0
M1718 793 541 163 163 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=98720 $D=0
M1719 794 542 164 164 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=103350 $D=0
M1720 645 647 793 163 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=98720 $D=0
M1721 646 648 794 164 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=103350 $D=0
M1722 647 635 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=99080 $D=0
M1723 648 636 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=103710 $D=0
M1724 649 645 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=99080 $D=0
M1725 650 646 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=103710 $D=0
M1726 163 643 649 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=99080 $D=0
M1727 164 644 650 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=103710 $D=0
M1728 652 157 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=99080 $D=0
M1729 653 651 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=103710 $D=0
M1730 651 649 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=99080 $D=0
M1731 158 650 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=103710 $D=0
M1732 163 652 651 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=99080 $D=0
M1733 164 653 158 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=103710 $D=0
M1734 655 654 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=99080 $D=0
M1735 656 159 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=103710 $D=0
M1736 163 659 657 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=99080 $D=0
M1737 164 660 658 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=103710 $D=0
M1738 661 115 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=99080 $D=0
M1739 662 116 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=103710 $D=0
M1740 659 115 654 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=99080 $D=0
M1741 660 116 159 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=103710 $D=0
M1742 655 661 659 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=99080 $D=0
M1743 656 662 660 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=103710 $D=0
M1744 663 657 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=99080 $D=0
M1745 664 658 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=103710 $D=0
M1746 160 657 5 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=99080 $D=0
M1747 654 658 6 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=103710 $D=0
M1748 115 663 160 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=99080 $D=0
M1749 116 664 654 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=103710 $D=0
M1750 665 160 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=99080 $D=0
M1751 666 654 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=103710 $D=0
M1752 667 657 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=99080 $D=0
M1753 668 658 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=103710 $D=0
M1754 203 657 665 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=99080 $D=0
M1755 204 658 666 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=103710 $D=0
M1756 5 667 203 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=99080 $D=0
M1757 6 668 204 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=103710 $D=0
M1758 669 161 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=99080 $D=0
M1759 670 161 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=103710 $D=0
M1760 671 161 203 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=99080 $D=0
M1761 672 161 204 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=103710 $D=0
M1762 12 669 671 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=99080 $D=0
M1763 13 670 672 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=103710 $D=0
M1764 673 162 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=99080 $D=0
M1765 674 162 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=103710 $D=0
M1766 162 162 671 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=99080 $D=0
M1767 162 162 672 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=103710 $D=0
M1768 5 673 162 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=99080 $D=0
M1769 6 674 162 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=103710 $D=0
M1770 675 111 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=99080 $D=0
M1771 676 111 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=103710 $D=0
M1772 163 675 677 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=99080 $D=0
M1773 164 676 678 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=103710 $D=0
M1774 679 111 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=99080 $D=0
M1775 680 111 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=103710 $D=0
M1776 681 677 162 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=99080 $D=0
M1777 682 678 162 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=103710 $D=0
M1778 163 681 781 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=99080 $D=0
M1779 164 682 782 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=103710 $D=0
M1780 683 781 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=99080 $D=0
M1781 684 782 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=103710 $D=0
M1782 681 675 683 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=99080 $D=0
M1783 682 676 684 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=103710 $D=0
M1784 685 679 683 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=99080 $D=0
M1785 686 680 684 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=103710 $D=0
M1786 163 689 687 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=99080 $D=0
M1787 164 690 688 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=103710 $D=0
M1788 689 111 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=99080 $D=0
M1789 690 111 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=103710 $D=0
M1790 783 685 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=99080 $D=0
M1791 784 686 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=103710 $D=0
M1792 691 689 783 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=99080 $D=0
M1793 692 690 784 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=103710 $D=0
M1794 163 691 115 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=99080 $D=0
M1795 164 692 116 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=103710 $D=0
M1796 785 115 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=99080 $D=0
M1797 786 116 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=103710 $D=0
M1798 691 687 785 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=99080 $D=0
M1799 692 688 786 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=103710 $D=0
.ENDS
***************************************
.SUBCKT ICV_29 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163
** N=805 EP=163 IP=1514 FDC=1800
M0 175 1 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=88570 $D=1
M1 176 1 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=93200 $D=1
M2 177 175 2 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=88570 $D=1
M3 178 176 3 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=93200 $D=1
M4 5 1 177 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=88570 $D=1
M5 6 1 178 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=93200 $D=1
M6 179 175 4 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=88570 $D=1
M7 180 176 4 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=93200 $D=1
M8 2 1 179 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=88570 $D=1
M9 3 1 180 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=93200 $D=1
M10 181 175 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=88570 $D=1
M11 182 176 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=93200 $D=1
M12 2 1 181 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=88570 $D=1
M13 3 1 182 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=93200 $D=1
M14 185 183 181 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=88570 $D=1
M15 186 184 182 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=93200 $D=1
M16 183 7 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=88570 $D=1
M17 184 7 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=93200 $D=1
M18 187 183 179 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=88570 $D=1
M19 188 184 180 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=93200 $D=1
M20 177 7 187 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=88570 $D=1
M21 178 7 188 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=93200 $D=1
M22 189 8 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=88570 $D=1
M23 190 8 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=93200 $D=1
M24 191 189 187 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=88570 $D=1
M25 192 190 188 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=93200 $D=1
M26 185 8 191 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=88570 $D=1
M27 186 8 192 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=93200 $D=1
M28 193 9 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=88570 $D=1
M29 194 9 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=93200 $D=1
M30 195 193 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=88570 $D=1
M31 196 194 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=93200 $D=1
M32 10 9 195 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=88570 $D=1
M33 11 9 196 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=93200 $D=1
M34 197 193 12 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=88570 $D=1
M35 198 194 13 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=93200 $D=1
M36 199 9 197 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=88570 $D=1
M37 200 9 198 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=93200 $D=1
M38 203 193 201 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=88570 $D=1
M39 204 194 202 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=93200 $D=1
M40 191 9 203 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=88570 $D=1
M41 192 9 204 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=93200 $D=1
M42 207 205 203 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=88570 $D=1
M43 208 206 204 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=93200 $D=1
M44 205 14 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=88570 $D=1
M45 206 14 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=93200 $D=1
M46 209 205 197 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=88570 $D=1
M47 210 206 198 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=93200 $D=1
M48 195 14 209 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=88570 $D=1
M49 196 14 210 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=93200 $D=1
M50 211 15 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=88570 $D=1
M51 212 15 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=93200 $D=1
M52 213 211 209 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=88570 $D=1
M53 214 212 210 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=93200 $D=1
M54 207 15 213 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=88570 $D=1
M55 208 15 214 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=93200 $D=1
M56 5 16 215 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=88570 $D=1
M57 6 16 216 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=93200 $D=1
M58 217 17 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=88570 $D=1
M59 218 17 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=93200 $D=1
M60 219 16 213 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=88570 $D=1
M61 220 16 214 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=93200 $D=1
M62 5 219 693 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=88570 $D=1
M63 6 220 694 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=93200 $D=1
M64 221 693 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=88570 $D=1
M65 222 694 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=93200 $D=1
M66 219 215 221 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=88570 $D=1
M67 220 216 222 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=93200 $D=1
M68 221 17 223 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=88570 $D=1
M69 222 17 224 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=93200 $D=1
M70 227 18 221 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=88570 $D=1
M71 228 18 222 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=93200 $D=1
M72 225 18 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=88570 $D=1
M73 226 18 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=93200 $D=1
M74 5 19 229 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=88570 $D=1
M75 6 19 230 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=93200 $D=1
M76 231 20 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=88570 $D=1
M77 232 20 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=93200 $D=1
M78 233 19 213 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=88570 $D=1
M79 234 19 214 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=93200 $D=1
M80 5 233 695 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=88570 $D=1
M81 6 234 696 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=93200 $D=1
M82 235 695 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=88570 $D=1
M83 236 696 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=93200 $D=1
M84 233 229 235 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=88570 $D=1
M85 234 230 236 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=93200 $D=1
M86 235 20 223 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=88570 $D=1
M87 236 20 224 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=93200 $D=1
M88 227 21 235 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=88570 $D=1
M89 228 21 236 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=93200 $D=1
M90 237 21 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=88570 $D=1
M91 238 21 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=93200 $D=1
M92 5 22 239 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=88570 $D=1
M93 6 22 240 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=93200 $D=1
M94 241 23 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=88570 $D=1
M95 242 23 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=93200 $D=1
M96 243 22 213 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=88570 $D=1
M97 244 22 214 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=93200 $D=1
M98 5 243 697 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=88570 $D=1
M99 6 244 698 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=93200 $D=1
M100 245 697 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=88570 $D=1
M101 246 698 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=93200 $D=1
M102 243 239 245 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=88570 $D=1
M103 244 240 246 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=93200 $D=1
M104 245 23 223 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=88570 $D=1
M105 246 23 224 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=93200 $D=1
M106 227 24 245 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=88570 $D=1
M107 228 24 246 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=93200 $D=1
M108 247 24 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=88570 $D=1
M109 248 24 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=93200 $D=1
M110 5 25 249 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=88570 $D=1
M111 6 25 250 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=93200 $D=1
M112 251 26 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=88570 $D=1
M113 252 26 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=93200 $D=1
M114 253 25 213 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=88570 $D=1
M115 254 25 214 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=93200 $D=1
M116 5 253 699 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=88570 $D=1
M117 6 254 700 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=93200 $D=1
M118 255 699 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=88570 $D=1
M119 256 700 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=93200 $D=1
M120 253 249 255 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=88570 $D=1
M121 254 250 256 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=93200 $D=1
M122 255 26 223 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=88570 $D=1
M123 256 26 224 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=93200 $D=1
M124 227 27 255 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=88570 $D=1
M125 228 27 256 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=93200 $D=1
M126 257 27 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=88570 $D=1
M127 258 27 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=93200 $D=1
M128 5 28 259 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=88570 $D=1
M129 6 28 260 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=93200 $D=1
M130 261 29 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=88570 $D=1
M131 262 29 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=93200 $D=1
M132 263 28 213 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=88570 $D=1
M133 264 28 214 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=93200 $D=1
M134 5 263 701 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=88570 $D=1
M135 6 264 702 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=93200 $D=1
M136 265 701 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=88570 $D=1
M137 266 702 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=93200 $D=1
M138 263 259 265 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=88570 $D=1
M139 264 260 266 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=93200 $D=1
M140 265 29 223 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=88570 $D=1
M141 266 29 224 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=93200 $D=1
M142 227 30 265 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=88570 $D=1
M143 228 30 266 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=93200 $D=1
M144 267 30 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=88570 $D=1
M145 268 30 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=93200 $D=1
M146 5 31 269 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=88570 $D=1
M147 6 31 270 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=93200 $D=1
M148 271 32 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=88570 $D=1
M149 272 32 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=93200 $D=1
M150 273 31 213 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=88570 $D=1
M151 274 31 214 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=93200 $D=1
M152 5 273 703 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=88570 $D=1
M153 6 274 704 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=93200 $D=1
M154 275 703 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=88570 $D=1
M155 276 704 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=93200 $D=1
M156 273 269 275 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=88570 $D=1
M157 274 270 276 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=93200 $D=1
M158 275 32 223 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=88570 $D=1
M159 276 32 224 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=93200 $D=1
M160 227 33 275 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=88570 $D=1
M161 228 33 276 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=93200 $D=1
M162 277 33 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=88570 $D=1
M163 278 33 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=93200 $D=1
M164 5 34 279 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=88570 $D=1
M165 6 34 280 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=93200 $D=1
M166 281 35 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=88570 $D=1
M167 282 35 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=93200 $D=1
M168 283 34 213 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=88570 $D=1
M169 284 34 214 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=93200 $D=1
M170 5 283 705 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=88570 $D=1
M171 6 284 706 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=93200 $D=1
M172 285 705 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=88570 $D=1
M173 286 706 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=93200 $D=1
M174 283 279 285 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=88570 $D=1
M175 284 280 286 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=93200 $D=1
M176 285 35 223 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=88570 $D=1
M177 286 35 224 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=93200 $D=1
M178 227 36 285 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=88570 $D=1
M179 228 36 286 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=93200 $D=1
M180 287 36 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=88570 $D=1
M181 288 36 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=93200 $D=1
M182 5 37 289 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=88570 $D=1
M183 6 37 290 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=93200 $D=1
M184 291 38 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=88570 $D=1
M185 292 38 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=93200 $D=1
M186 293 37 213 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=88570 $D=1
M187 294 37 214 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=93200 $D=1
M188 5 293 707 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=88570 $D=1
M189 6 294 708 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=93200 $D=1
M190 295 707 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=88570 $D=1
M191 296 708 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=93200 $D=1
M192 293 289 295 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=88570 $D=1
M193 294 290 296 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=93200 $D=1
M194 295 38 223 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=88570 $D=1
M195 296 38 224 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=93200 $D=1
M196 227 39 295 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=88570 $D=1
M197 228 39 296 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=93200 $D=1
M198 297 39 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=88570 $D=1
M199 298 39 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=93200 $D=1
M200 5 40 299 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=88570 $D=1
M201 6 40 300 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=93200 $D=1
M202 301 41 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=88570 $D=1
M203 302 41 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=93200 $D=1
M204 303 40 213 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=88570 $D=1
M205 304 40 214 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=93200 $D=1
M206 5 303 709 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=88570 $D=1
M207 6 304 710 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=93200 $D=1
M208 305 709 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=88570 $D=1
M209 306 710 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=93200 $D=1
M210 303 299 305 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=88570 $D=1
M211 304 300 306 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=93200 $D=1
M212 305 41 223 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=88570 $D=1
M213 306 41 224 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=93200 $D=1
M214 227 42 305 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=88570 $D=1
M215 228 42 306 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=93200 $D=1
M216 307 42 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=88570 $D=1
M217 308 42 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=93200 $D=1
M218 5 43 309 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=88570 $D=1
M219 6 43 310 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=93200 $D=1
M220 311 44 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=88570 $D=1
M221 312 44 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=93200 $D=1
M222 313 43 213 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=88570 $D=1
M223 314 43 214 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=93200 $D=1
M224 5 313 711 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=88570 $D=1
M225 6 314 712 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=93200 $D=1
M226 315 711 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=88570 $D=1
M227 316 712 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=93200 $D=1
M228 313 309 315 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=88570 $D=1
M229 314 310 316 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=93200 $D=1
M230 315 44 223 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=88570 $D=1
M231 316 44 224 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=93200 $D=1
M232 227 45 315 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=88570 $D=1
M233 228 45 316 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=93200 $D=1
M234 317 45 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=88570 $D=1
M235 318 45 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=93200 $D=1
M236 5 46 319 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=88570 $D=1
M237 6 46 320 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=93200 $D=1
M238 321 47 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=88570 $D=1
M239 322 47 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=93200 $D=1
M240 323 46 213 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=88570 $D=1
M241 324 46 214 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=93200 $D=1
M242 5 323 713 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=88570 $D=1
M243 6 324 714 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=93200 $D=1
M244 325 713 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=88570 $D=1
M245 326 714 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=93200 $D=1
M246 323 319 325 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=88570 $D=1
M247 324 320 326 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=93200 $D=1
M248 325 47 223 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=88570 $D=1
M249 326 47 224 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=93200 $D=1
M250 227 48 325 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=88570 $D=1
M251 228 48 326 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=93200 $D=1
M252 327 48 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=88570 $D=1
M253 328 48 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=93200 $D=1
M254 5 49 329 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=88570 $D=1
M255 6 49 330 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=93200 $D=1
M256 331 50 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=88570 $D=1
M257 332 50 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=93200 $D=1
M258 333 49 213 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=88570 $D=1
M259 334 49 214 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=93200 $D=1
M260 5 333 715 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=88570 $D=1
M261 6 334 716 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=93200 $D=1
M262 335 715 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=88570 $D=1
M263 336 716 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=93200 $D=1
M264 333 329 335 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=88570 $D=1
M265 334 330 336 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=93200 $D=1
M266 335 50 223 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=88570 $D=1
M267 336 50 224 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=93200 $D=1
M268 227 51 335 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=88570 $D=1
M269 228 51 336 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=93200 $D=1
M270 337 51 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=88570 $D=1
M271 338 51 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=93200 $D=1
M272 5 52 339 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=88570 $D=1
M273 6 52 340 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=93200 $D=1
M274 341 53 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=88570 $D=1
M275 342 53 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=93200 $D=1
M276 343 52 213 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=88570 $D=1
M277 344 52 214 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=93200 $D=1
M278 5 343 717 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=88570 $D=1
M279 6 344 718 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=93200 $D=1
M280 345 717 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=88570 $D=1
M281 346 718 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=93200 $D=1
M282 343 339 345 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=88570 $D=1
M283 344 340 346 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=93200 $D=1
M284 345 53 223 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=88570 $D=1
M285 346 53 224 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=93200 $D=1
M286 227 54 345 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=88570 $D=1
M287 228 54 346 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=93200 $D=1
M288 347 54 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=88570 $D=1
M289 348 54 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=93200 $D=1
M290 5 55 349 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=88570 $D=1
M291 6 55 350 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=93200 $D=1
M292 351 56 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=88570 $D=1
M293 352 56 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=93200 $D=1
M294 353 55 213 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=88570 $D=1
M295 354 55 214 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=93200 $D=1
M296 5 353 719 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=88570 $D=1
M297 6 354 720 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=93200 $D=1
M298 355 719 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=88570 $D=1
M299 356 720 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=93200 $D=1
M300 353 349 355 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=88570 $D=1
M301 354 350 356 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=93200 $D=1
M302 355 56 223 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=88570 $D=1
M303 356 56 224 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=93200 $D=1
M304 227 57 355 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=88570 $D=1
M305 228 57 356 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=93200 $D=1
M306 357 57 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=88570 $D=1
M307 358 57 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=93200 $D=1
M308 5 58 359 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=88570 $D=1
M309 6 58 360 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=93200 $D=1
M310 361 59 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=88570 $D=1
M311 362 59 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=93200 $D=1
M312 363 58 213 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=88570 $D=1
M313 364 58 214 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=93200 $D=1
M314 5 363 721 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=88570 $D=1
M315 6 364 722 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=93200 $D=1
M316 365 721 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=88570 $D=1
M317 366 722 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=93200 $D=1
M318 363 359 365 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=88570 $D=1
M319 364 360 366 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=93200 $D=1
M320 365 59 223 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=88570 $D=1
M321 366 59 224 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=93200 $D=1
M322 227 60 365 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=88570 $D=1
M323 228 60 366 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=93200 $D=1
M324 367 60 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=88570 $D=1
M325 368 60 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=93200 $D=1
M326 5 61 369 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=88570 $D=1
M327 6 61 370 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=93200 $D=1
M328 371 62 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=88570 $D=1
M329 372 62 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=93200 $D=1
M330 373 61 213 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=88570 $D=1
M331 374 61 214 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=93200 $D=1
M332 5 373 723 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=88570 $D=1
M333 6 374 724 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=93200 $D=1
M334 375 723 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=88570 $D=1
M335 376 724 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=93200 $D=1
M336 373 369 375 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=88570 $D=1
M337 374 370 376 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=93200 $D=1
M338 375 62 223 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=88570 $D=1
M339 376 62 224 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=93200 $D=1
M340 227 63 375 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=88570 $D=1
M341 228 63 376 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=93200 $D=1
M342 377 63 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=88570 $D=1
M343 378 63 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=93200 $D=1
M344 5 64 379 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=88570 $D=1
M345 6 64 380 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=93200 $D=1
M346 381 65 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=88570 $D=1
M347 382 65 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=93200 $D=1
M348 383 64 213 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=88570 $D=1
M349 384 64 214 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=93200 $D=1
M350 5 383 725 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=88570 $D=1
M351 6 384 726 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=93200 $D=1
M352 385 725 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=88570 $D=1
M353 386 726 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=93200 $D=1
M354 383 379 385 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=88570 $D=1
M355 384 380 386 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=93200 $D=1
M356 385 65 223 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=88570 $D=1
M357 386 65 224 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=93200 $D=1
M358 227 66 385 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=88570 $D=1
M359 228 66 386 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=93200 $D=1
M360 387 66 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=88570 $D=1
M361 388 66 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=93200 $D=1
M362 5 67 389 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=88570 $D=1
M363 6 67 390 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=93200 $D=1
M364 391 68 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=88570 $D=1
M365 392 68 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=93200 $D=1
M366 393 67 213 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=88570 $D=1
M367 394 67 214 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=93200 $D=1
M368 5 393 727 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=88570 $D=1
M369 6 394 728 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=93200 $D=1
M370 395 727 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=88570 $D=1
M371 396 728 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=93200 $D=1
M372 393 389 395 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=88570 $D=1
M373 394 390 396 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=93200 $D=1
M374 395 68 223 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=88570 $D=1
M375 396 68 224 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=93200 $D=1
M376 227 69 395 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=88570 $D=1
M377 228 69 396 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=93200 $D=1
M378 397 69 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=88570 $D=1
M379 398 69 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=93200 $D=1
M380 5 70 399 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=88570 $D=1
M381 6 70 400 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=93200 $D=1
M382 401 71 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=88570 $D=1
M383 402 71 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=93200 $D=1
M384 403 70 213 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=88570 $D=1
M385 404 70 214 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=93200 $D=1
M386 5 403 729 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=88570 $D=1
M387 6 404 730 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=93200 $D=1
M388 405 729 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=88570 $D=1
M389 406 730 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=93200 $D=1
M390 403 399 405 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=88570 $D=1
M391 404 400 406 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=93200 $D=1
M392 405 71 223 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=88570 $D=1
M393 406 71 224 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=93200 $D=1
M394 227 72 405 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=88570 $D=1
M395 228 72 406 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=93200 $D=1
M396 407 72 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=88570 $D=1
M397 408 72 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=93200 $D=1
M398 5 73 409 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=88570 $D=1
M399 6 73 410 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=93200 $D=1
M400 411 74 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=88570 $D=1
M401 412 74 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=93200 $D=1
M402 413 73 213 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=88570 $D=1
M403 414 73 214 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=93200 $D=1
M404 5 413 731 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=88570 $D=1
M405 6 414 732 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=93200 $D=1
M406 415 731 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=88570 $D=1
M407 416 732 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=93200 $D=1
M408 413 409 415 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=88570 $D=1
M409 414 410 416 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=93200 $D=1
M410 415 74 223 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=88570 $D=1
M411 416 74 224 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=93200 $D=1
M412 227 75 415 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=88570 $D=1
M413 228 75 416 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=93200 $D=1
M414 417 75 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=88570 $D=1
M415 418 75 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=93200 $D=1
M416 5 76 419 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=88570 $D=1
M417 6 76 420 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=93200 $D=1
M418 421 77 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=88570 $D=1
M419 422 77 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=93200 $D=1
M420 423 76 213 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=88570 $D=1
M421 424 76 214 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=93200 $D=1
M422 5 423 733 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=88570 $D=1
M423 6 424 734 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=93200 $D=1
M424 425 733 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=88570 $D=1
M425 426 734 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=93200 $D=1
M426 423 419 425 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=88570 $D=1
M427 424 420 426 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=93200 $D=1
M428 425 77 223 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=88570 $D=1
M429 426 77 224 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=93200 $D=1
M430 227 78 425 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=88570 $D=1
M431 228 78 426 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=93200 $D=1
M432 427 78 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=88570 $D=1
M433 428 78 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=93200 $D=1
M434 5 79 429 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=88570 $D=1
M435 6 79 430 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=93200 $D=1
M436 431 80 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=88570 $D=1
M437 432 80 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=93200 $D=1
M438 433 79 213 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=88570 $D=1
M439 434 79 214 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=93200 $D=1
M440 5 433 735 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=88570 $D=1
M441 6 434 736 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=93200 $D=1
M442 435 735 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=88570 $D=1
M443 436 736 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=93200 $D=1
M444 433 429 435 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=88570 $D=1
M445 434 430 436 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=93200 $D=1
M446 435 80 223 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=88570 $D=1
M447 436 80 224 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=93200 $D=1
M448 227 81 435 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=88570 $D=1
M449 228 81 436 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=93200 $D=1
M450 437 81 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=88570 $D=1
M451 438 81 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=93200 $D=1
M452 5 82 439 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=88570 $D=1
M453 6 82 440 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=93200 $D=1
M454 441 83 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=88570 $D=1
M455 442 83 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=93200 $D=1
M456 443 82 213 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=88570 $D=1
M457 444 82 214 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=93200 $D=1
M458 5 443 737 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=88570 $D=1
M459 6 444 738 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=93200 $D=1
M460 445 737 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=88570 $D=1
M461 446 738 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=93200 $D=1
M462 443 439 445 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=88570 $D=1
M463 444 440 446 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=93200 $D=1
M464 445 83 223 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=88570 $D=1
M465 446 83 224 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=93200 $D=1
M466 227 84 445 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=88570 $D=1
M467 228 84 446 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=93200 $D=1
M468 447 84 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=88570 $D=1
M469 448 84 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=93200 $D=1
M470 5 85 449 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=88570 $D=1
M471 6 85 450 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=93200 $D=1
M472 451 86 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=88570 $D=1
M473 452 86 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=93200 $D=1
M474 453 85 213 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=88570 $D=1
M475 454 85 214 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=93200 $D=1
M476 5 453 739 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=88570 $D=1
M477 6 454 740 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=93200 $D=1
M478 455 739 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=88570 $D=1
M479 456 740 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=93200 $D=1
M480 453 449 455 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=88570 $D=1
M481 454 450 456 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=93200 $D=1
M482 455 86 223 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=88570 $D=1
M483 456 86 224 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=93200 $D=1
M484 227 87 455 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=88570 $D=1
M485 228 87 456 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=93200 $D=1
M486 457 87 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=88570 $D=1
M487 458 87 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=93200 $D=1
M488 5 88 459 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=88570 $D=1
M489 6 88 460 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=93200 $D=1
M490 461 89 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=88570 $D=1
M491 462 89 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=93200 $D=1
M492 463 88 213 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=88570 $D=1
M493 464 88 214 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=93200 $D=1
M494 5 463 741 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=88570 $D=1
M495 6 464 742 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=93200 $D=1
M496 465 741 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=88570 $D=1
M497 466 742 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=93200 $D=1
M498 463 459 465 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=88570 $D=1
M499 464 460 466 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=93200 $D=1
M500 465 89 223 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=88570 $D=1
M501 466 89 224 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=93200 $D=1
M502 227 90 465 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=88570 $D=1
M503 228 90 466 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=93200 $D=1
M504 467 90 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=88570 $D=1
M505 468 90 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=93200 $D=1
M506 5 91 469 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=88570 $D=1
M507 6 91 470 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=93200 $D=1
M508 471 92 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=88570 $D=1
M509 472 92 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=93200 $D=1
M510 473 91 213 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=88570 $D=1
M511 474 91 214 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=93200 $D=1
M512 5 473 743 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=88570 $D=1
M513 6 474 744 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=93200 $D=1
M514 475 743 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=88570 $D=1
M515 476 744 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=93200 $D=1
M516 473 469 475 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=88570 $D=1
M517 474 470 476 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=93200 $D=1
M518 475 92 223 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=88570 $D=1
M519 476 92 224 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=93200 $D=1
M520 227 93 475 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=88570 $D=1
M521 228 93 476 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=93200 $D=1
M522 477 93 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=88570 $D=1
M523 478 93 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=93200 $D=1
M524 5 94 479 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=88570 $D=1
M525 6 94 480 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=93200 $D=1
M526 481 95 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=88570 $D=1
M527 482 95 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=93200 $D=1
M528 483 94 213 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=88570 $D=1
M529 484 94 214 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=93200 $D=1
M530 5 483 745 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=88570 $D=1
M531 6 484 746 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=93200 $D=1
M532 485 745 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=88570 $D=1
M533 486 746 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=93200 $D=1
M534 483 479 485 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=88570 $D=1
M535 484 480 486 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=93200 $D=1
M536 485 95 223 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=88570 $D=1
M537 486 95 224 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=93200 $D=1
M538 227 96 485 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=88570 $D=1
M539 228 96 486 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=93200 $D=1
M540 487 96 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=88570 $D=1
M541 488 96 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=93200 $D=1
M542 5 97 489 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=88570 $D=1
M543 6 97 490 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=93200 $D=1
M544 491 98 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=88570 $D=1
M545 492 98 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=93200 $D=1
M546 493 97 213 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=88570 $D=1
M547 494 97 214 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=93200 $D=1
M548 5 493 747 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=88570 $D=1
M549 6 494 748 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=93200 $D=1
M550 495 747 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=88570 $D=1
M551 496 748 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=93200 $D=1
M552 493 489 495 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=88570 $D=1
M553 494 490 496 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=93200 $D=1
M554 495 98 223 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=88570 $D=1
M555 496 98 224 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=93200 $D=1
M556 227 99 495 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=88570 $D=1
M557 228 99 496 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=93200 $D=1
M558 497 99 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=88570 $D=1
M559 498 99 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=93200 $D=1
M560 5 100 499 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=88570 $D=1
M561 6 100 500 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=93200 $D=1
M562 501 101 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=88570 $D=1
M563 502 101 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=93200 $D=1
M564 503 100 213 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=88570 $D=1
M565 504 100 214 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=93200 $D=1
M566 5 503 749 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=88570 $D=1
M567 6 504 750 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=93200 $D=1
M568 505 749 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=88570 $D=1
M569 506 750 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=93200 $D=1
M570 503 499 505 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=88570 $D=1
M571 504 500 506 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=93200 $D=1
M572 505 101 223 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=88570 $D=1
M573 506 101 224 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=93200 $D=1
M574 227 102 505 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=88570 $D=1
M575 228 102 506 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=93200 $D=1
M576 507 102 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=88570 $D=1
M577 508 102 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=93200 $D=1
M578 5 103 509 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=88570 $D=1
M579 6 103 510 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=93200 $D=1
M580 511 104 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=88570 $D=1
M581 512 104 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=93200 $D=1
M582 513 103 213 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=88570 $D=1
M583 514 103 214 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=93200 $D=1
M584 5 513 751 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=88570 $D=1
M585 6 514 752 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=93200 $D=1
M586 515 751 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=88570 $D=1
M587 516 752 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=93200 $D=1
M588 513 509 515 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=88570 $D=1
M589 514 510 516 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=93200 $D=1
M590 515 104 223 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=88570 $D=1
M591 516 104 224 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=93200 $D=1
M592 227 105 515 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=88570 $D=1
M593 228 105 516 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=93200 $D=1
M594 517 105 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=88570 $D=1
M595 518 105 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=93200 $D=1
M596 5 106 519 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=88570 $D=1
M597 6 106 520 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=93200 $D=1
M598 521 107 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=88570 $D=1
M599 522 107 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=93200 $D=1
M600 523 106 213 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=88570 $D=1
M601 524 106 214 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=93200 $D=1
M602 5 523 753 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=88570 $D=1
M603 6 524 754 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=93200 $D=1
M604 525 753 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=88570 $D=1
M605 526 754 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=93200 $D=1
M606 523 519 525 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=88570 $D=1
M607 524 520 526 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=93200 $D=1
M608 525 107 223 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=88570 $D=1
M609 526 107 224 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=93200 $D=1
M610 227 108 525 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=88570 $D=1
M611 228 108 526 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=93200 $D=1
M612 527 108 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=88570 $D=1
M613 528 108 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=93200 $D=1
M614 5 109 529 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=88570 $D=1
M615 6 109 530 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=93200 $D=1
M616 531 110 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=88570 $D=1
M617 532 110 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=93200 $D=1
M618 5 110 223 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=88570 $D=1
M619 6 110 224 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=93200 $D=1
M620 227 109 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=88570 $D=1
M621 228 109 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=93200 $D=1
M622 5 535 533 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=88570 $D=1
M623 6 536 534 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=93200 $D=1
M624 535 111 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=88570 $D=1
M625 536 111 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=93200 $D=1
M626 755 223 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=88570 $D=1
M627 756 224 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=93200 $D=1
M628 537 533 755 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=88570 $D=1
M629 538 534 756 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=93200 $D=1
M630 5 537 539 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=88570 $D=1
M631 6 538 540 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=93200 $D=1
M632 757 539 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=88570 $D=1
M633 758 540 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=93200 $D=1
M634 537 535 757 5 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=88570 $D=1
M635 538 536 758 6 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=93200 $D=1
M636 5 543 541 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=88570 $D=1
M637 6 544 542 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=93200 $D=1
M638 543 111 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=88570 $D=1
M639 544 111 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=93200 $D=1
M640 759 227 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=88570 $D=1
M641 760 228 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=93200 $D=1
M642 545 541 759 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=88570 $D=1
M643 546 542 760 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=93200 $D=1
M644 5 545 112 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=88570 $D=1
M645 6 546 113 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=93200 $D=1
M646 761 112 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=88570 $D=1
M647 762 113 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=93200 $D=1
M648 545 543 761 5 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=88570 $D=1
M649 546 544 762 6 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=93200 $D=1
M650 547 114 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=88570 $D=1
M651 548 114 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=93200 $D=1
M652 549 547 539 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=88570 $D=1
M653 550 548 540 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=93200 $D=1
M654 115 114 549 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=88570 $D=1
M655 116 114 550 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=93200 $D=1
M656 551 117 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=88570 $D=1
M657 552 117 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=93200 $D=1
M658 553 551 112 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=88570 $D=1
M659 554 552 113 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=93200 $D=1
M660 763 117 553 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=88570 $D=1
M661 764 117 554 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=93200 $D=1
M662 5 112 763 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=88570 $D=1
M663 6 113 764 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=93200 $D=1
M664 555 118 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=88570 $D=1
M665 556 118 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=93200 $D=1
M666 557 555 553 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=88570 $D=1
M667 558 556 554 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=93200 $D=1
M668 10 118 557 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=88570 $D=1
M669 11 118 558 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=93200 $D=1
M670 560 559 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=88570 $D=1
M671 561 119 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=93200 $D=1
M672 5 564 562 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=88570 $D=1
M673 6 565 563 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=93200 $D=1
M674 566 549 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=88570 $D=1
M675 567 550 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=93200 $D=1
M676 564 566 559 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=88570 $D=1
M677 565 567 119 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=93200 $D=1
M678 560 549 564 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=88570 $D=1
M679 561 550 565 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=93200 $D=1
M680 568 562 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=88570 $D=1
M681 569 563 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=93200 $D=1
M682 570 568 557 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=88570 $D=1
M683 559 569 558 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=93200 $D=1
M684 549 562 570 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=88570 $D=1
M685 550 563 559 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=93200 $D=1
M686 571 570 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=88570 $D=1
M687 572 559 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=93200 $D=1
M688 573 562 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=88570 $D=1
M689 574 563 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=93200 $D=1
M690 575 573 571 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=88570 $D=1
M691 576 574 572 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=93200 $D=1
M692 557 562 575 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=88570 $D=1
M693 558 563 576 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=93200 $D=1
M694 577 549 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=88570 $D=1
M695 578 550 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=93200 $D=1
M696 5 557 577 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=88570 $D=1
M697 6 558 578 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=93200 $D=1
M698 579 575 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=88570 $D=1
M699 580 576 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=93200 $D=1
M700 794 549 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=88570 $D=1
M701 795 550 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=93200 $D=1
M702 581 557 794 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=88570 $D=1
M703 582 558 795 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=93200 $D=1
M704 796 549 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=88570 $D=1
M705 797 550 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=93200 $D=1
M706 583 557 796 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=88570 $D=1
M707 584 558 797 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=93200 $D=1
M708 587 549 585 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=88570 $D=1
M709 588 550 586 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=93200 $D=1
M710 585 557 587 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=88570 $D=1
M711 586 558 588 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=93200 $D=1
M712 5 583 585 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=88570 $D=1
M713 6 584 586 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=93200 $D=1
M714 589 121 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=88570 $D=1
M715 590 121 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=93200 $D=1
M716 591 589 577 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=88570 $D=1
M717 592 590 578 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=93200 $D=1
M718 581 121 591 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=88570 $D=1
M719 582 121 592 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=93200 $D=1
M720 593 589 579 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=88570 $D=1
M721 594 590 580 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=93200 $D=1
M722 587 121 593 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=88570 $D=1
M723 588 121 594 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=93200 $D=1
M724 595 122 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=88570 $D=1
M725 596 122 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=93200 $D=1
M726 597 595 593 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=88570 $D=1
M727 598 596 594 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=93200 $D=1
M728 591 122 597 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=88570 $D=1
M729 592 122 598 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=93200 $D=1
M730 12 597 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=88570 $D=1
M731 13 598 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=93200 $D=1
M732 599 123 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=88570 $D=1
M733 600 123 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=93200 $D=1
M734 601 599 124 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=88570 $D=1
M735 602 600 125 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=93200 $D=1
M736 126 123 601 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=88570 $D=1
M737 127 123 602 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=93200 $D=1
M738 603 123 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=88570 $D=1
M739 604 123 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=93200 $D=1
M740 609 603 128 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=88570 $D=1
M741 610 604 130 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=93200 $D=1
M742 131 123 609 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=88570 $D=1
M743 129 123 610 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=93200 $D=1
M744 611 123 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=88570 $D=1
M745 612 123 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=93200 $D=1
M746 613 611 132 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=88570 $D=1
M747 614 612 133 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=93200 $D=1
M748 134 123 613 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=88570 $D=1
M749 135 123 614 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=93200 $D=1
M750 615 123 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=88570 $D=1
M751 616 123 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=93200 $D=1
M752 617 615 136 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=88570 $D=1
M753 618 616 137 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=93200 $D=1
M754 138 123 617 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=88570 $D=1
M755 139 123 618 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=93200 $D=1
M756 619 123 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=88570 $D=1
M757 620 123 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=93200 $D=1
M758 621 619 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=88570 $D=1
M759 622 620 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=93200 $D=1
M760 140 123 621 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=88570 $D=1
M761 141 123 622 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=93200 $D=1
M762 5 549 776 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=88570 $D=1
M763 6 550 777 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=93200 $D=1
M764 127 776 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=88570 $D=1
M765 124 777 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=93200 $D=1
M766 623 142 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=88570 $D=1
M767 624 142 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=93200 $D=1
M768 143 623 127 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=88570 $D=1
M769 144 624 124 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=93200 $D=1
M770 601 142 143 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=88570 $D=1
M771 602 142 144 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=93200 $D=1
M772 625 145 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=88570 $D=1
M773 626 145 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=93200 $D=1
M774 120 625 143 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=88570 $D=1
M775 146 626 144 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=93200 $D=1
M776 609 145 120 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=88570 $D=1
M777 610 145 146 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=93200 $D=1
M778 627 147 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=88570 $D=1
M779 628 147 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=93200 $D=1
M780 148 627 120 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=88570 $D=1
M781 149 628 146 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=93200 $D=1
M782 613 147 148 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=88570 $D=1
M783 614 147 149 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=93200 $D=1
M784 629 150 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=88570 $D=1
M785 630 150 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=93200 $D=1
M786 151 629 148 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=88570 $D=1
M787 152 630 149 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=93200 $D=1
M788 617 150 151 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=88570 $D=1
M789 618 150 152 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=93200 $D=1
M790 631 153 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=88570 $D=1
M791 632 153 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=93200 $D=1
M792 199 631 151 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=88570 $D=1
M793 200 632 152 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=93200 $D=1
M794 621 153 199 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=88570 $D=1
M795 622 153 200 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=93200 $D=1
M796 633 154 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=88570 $D=1
M797 634 154 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=93200 $D=1
M798 635 633 112 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=88570 $D=1
M799 636 634 113 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=93200 $D=1
M800 10 154 635 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=88570 $D=1
M801 11 154 636 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=93200 $D=1
M802 798 539 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=88570 $D=1
M803 799 540 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=93200 $D=1
M804 637 635 798 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=88570 $D=1
M805 638 636 799 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=93200 $D=1
M806 641 539 639 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=88570 $D=1
M807 642 540 640 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=93200 $D=1
M808 639 635 641 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=88570 $D=1
M809 640 636 642 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=93200 $D=1
M810 5 637 639 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=88570 $D=1
M811 6 638 640 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=93200 $D=1
M812 800 643 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=88570 $D=1
M813 801 644 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=93200 $D=1
M814 778 641 800 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=88570 $D=1
M815 779 642 801 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=93200 $D=1
M816 644 778 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=88570 $D=1
M817 155 779 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=93200 $D=1
M818 645 539 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=88570 $D=1
M819 646 540 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=93200 $D=1
M820 5 647 645 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=88570 $D=1
M821 6 648 646 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=93200 $D=1
M822 647 635 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=88570 $D=1
M823 648 636 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=93200 $D=1
M824 802 645 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=88570 $D=1
M825 803 646 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=93200 $D=1
M826 649 643 802 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=88570 $D=1
M827 650 644 803 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=93200 $D=1
M828 652 156 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=88570 $D=1
M829 653 651 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=93200 $D=1
M830 804 649 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=88570 $D=1
M831 805 650 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=93200 $D=1
M832 651 652 804 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=88570 $D=1
M833 157 653 805 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=93200 $D=1
M834 655 654 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=88570 $D=1
M835 656 158 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=93200 $D=1
M836 5 659 657 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=88570 $D=1
M837 6 660 658 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=93200 $D=1
M838 661 115 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=88570 $D=1
M839 662 116 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=93200 $D=1
M840 659 661 654 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=88570 $D=1
M841 660 662 158 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=93200 $D=1
M842 655 115 659 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=88570 $D=1
M843 656 116 660 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=93200 $D=1
M844 663 657 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=88570 $D=1
M845 664 658 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=93200 $D=1
M846 159 663 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=88570 $D=1
M847 654 664 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=93200 $D=1
M848 115 657 159 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=88570 $D=1
M849 116 658 654 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=93200 $D=1
M850 665 159 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=88570 $D=1
M851 666 654 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=93200 $D=1
M852 667 657 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=88570 $D=1
M853 668 658 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=93200 $D=1
M854 201 667 665 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=88570 $D=1
M855 202 668 666 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=93200 $D=1
M856 5 657 201 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=88570 $D=1
M857 6 658 202 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=93200 $D=1
M858 669 160 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=88570 $D=1
M859 670 160 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=93200 $D=1
M860 671 669 201 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=88570 $D=1
M861 672 670 202 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=93200 $D=1
M862 12 160 671 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=88570 $D=1
M863 13 160 672 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=93200 $D=1
M864 673 161 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=88570 $D=1
M865 674 161 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=93200 $D=1
M866 161 673 671 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=88570 $D=1
M867 161 674 672 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=93200 $D=1
M868 5 161 161 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=88570 $D=1
M869 6 161 161 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=93200 $D=1
M870 675 111 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=88570 $D=1
M871 676 111 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=93200 $D=1
M872 5 675 677 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=88570 $D=1
M873 6 676 678 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=93200 $D=1
M874 679 111 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=88570 $D=1
M875 680 111 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=93200 $D=1
M876 681 675 161 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=88570 $D=1
M877 682 676 161 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=93200 $D=1
M878 5 681 780 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=88570 $D=1
M879 6 682 781 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=93200 $D=1
M880 683 780 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=88570 $D=1
M881 684 781 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=93200 $D=1
M882 681 677 683 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=88570 $D=1
M883 682 678 684 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=93200 $D=1
M884 685 111 683 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=88570 $D=1
M885 686 111 684 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=93200 $D=1
M886 5 689 687 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=88570 $D=1
M887 6 690 688 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=93200 $D=1
M888 689 111 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=88570 $D=1
M889 690 111 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=93200 $D=1
M890 782 685 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=88570 $D=1
M891 783 686 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=93200 $D=1
M892 691 687 782 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=88570 $D=1
M893 692 688 783 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=93200 $D=1
M894 5 691 115 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=88570 $D=1
M895 6 692 116 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=93200 $D=1
M896 784 115 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=88570 $D=1
M897 785 116 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=93200 $D=1
M898 691 689 784 5 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=88570 $D=1
M899 692 690 785 6 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=93200 $D=1
M900 175 1 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=89820 $D=0
M901 176 1 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=94450 $D=0
M902 177 1 2 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=89820 $D=0
M903 178 1 3 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=94450 $D=0
M904 5 175 177 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=89820 $D=0
M905 6 176 178 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=94450 $D=0
M906 179 1 4 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=89820 $D=0
M907 180 1 4 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=94450 $D=0
M908 2 175 179 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=89820 $D=0
M909 3 176 180 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=94450 $D=0
M910 181 1 5 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=89820 $D=0
M911 182 1 6 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=94450 $D=0
M912 2 175 181 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=89820 $D=0
M913 3 176 182 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=94450 $D=0
M914 185 7 181 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=89820 $D=0
M915 186 7 182 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=94450 $D=0
M916 183 7 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=89820 $D=0
M917 184 7 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=94450 $D=0
M918 187 7 179 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=89820 $D=0
M919 188 7 180 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=94450 $D=0
M920 177 183 187 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=89820 $D=0
M921 178 184 188 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=94450 $D=0
M922 189 8 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=89820 $D=0
M923 190 8 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=94450 $D=0
M924 191 8 187 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=89820 $D=0
M925 192 8 188 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=94450 $D=0
M926 185 189 191 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=89820 $D=0
M927 186 190 192 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=94450 $D=0
M928 193 9 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=89820 $D=0
M929 194 9 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=94450 $D=0
M930 195 9 5 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=89820 $D=0
M931 196 9 6 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=94450 $D=0
M932 10 193 195 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=89820 $D=0
M933 11 194 196 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=94450 $D=0
M934 197 9 12 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=89820 $D=0
M935 198 9 13 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=94450 $D=0
M936 199 193 197 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=89820 $D=0
M937 200 194 198 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=94450 $D=0
M938 203 9 201 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=89820 $D=0
M939 204 9 202 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=94450 $D=0
M940 191 193 203 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=89820 $D=0
M941 192 194 204 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=94450 $D=0
M942 207 14 203 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=89820 $D=0
M943 208 14 204 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=94450 $D=0
M944 205 14 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=89820 $D=0
M945 206 14 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=94450 $D=0
M946 209 14 197 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=89820 $D=0
M947 210 14 198 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=94450 $D=0
M948 195 205 209 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=89820 $D=0
M949 196 206 210 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=94450 $D=0
M950 211 15 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=89820 $D=0
M951 212 15 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=94450 $D=0
M952 213 15 209 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=89820 $D=0
M953 214 15 210 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=94450 $D=0
M954 207 211 213 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=89820 $D=0
M955 208 212 214 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=94450 $D=0
M956 162 16 215 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=89820 $D=0
M957 163 16 216 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=94450 $D=0
M958 217 17 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=89820 $D=0
M959 218 17 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=94450 $D=0
M960 219 215 213 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=89820 $D=0
M961 220 216 214 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=94450 $D=0
M962 162 219 693 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=89820 $D=0
M963 163 220 694 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=94450 $D=0
M964 221 693 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=89820 $D=0
M965 222 694 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=94450 $D=0
M966 219 16 221 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=89820 $D=0
M967 220 16 222 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=94450 $D=0
M968 221 217 223 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=89820 $D=0
M969 222 218 224 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=94450 $D=0
M970 227 225 221 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=89820 $D=0
M971 228 226 222 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=94450 $D=0
M972 225 18 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=89820 $D=0
M973 226 18 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=94450 $D=0
M974 162 19 229 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=89820 $D=0
M975 163 19 230 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=94450 $D=0
M976 231 20 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=89820 $D=0
M977 232 20 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=94450 $D=0
M978 233 229 213 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=89820 $D=0
M979 234 230 214 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=94450 $D=0
M980 162 233 695 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=89820 $D=0
M981 163 234 696 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=94450 $D=0
M982 235 695 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=89820 $D=0
M983 236 696 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=94450 $D=0
M984 233 19 235 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=89820 $D=0
M985 234 19 236 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=94450 $D=0
M986 235 231 223 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=89820 $D=0
M987 236 232 224 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=94450 $D=0
M988 227 237 235 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=89820 $D=0
M989 228 238 236 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=94450 $D=0
M990 237 21 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=89820 $D=0
M991 238 21 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=94450 $D=0
M992 162 22 239 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=89820 $D=0
M993 163 22 240 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=94450 $D=0
M994 241 23 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=89820 $D=0
M995 242 23 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=94450 $D=0
M996 243 239 213 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=89820 $D=0
M997 244 240 214 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=94450 $D=0
M998 162 243 697 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=89820 $D=0
M999 163 244 698 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=94450 $D=0
M1000 245 697 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=89820 $D=0
M1001 246 698 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=94450 $D=0
M1002 243 22 245 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=89820 $D=0
M1003 244 22 246 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=94450 $D=0
M1004 245 241 223 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=89820 $D=0
M1005 246 242 224 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=94450 $D=0
M1006 227 247 245 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=89820 $D=0
M1007 228 248 246 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=94450 $D=0
M1008 247 24 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=89820 $D=0
M1009 248 24 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=94450 $D=0
M1010 162 25 249 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=89820 $D=0
M1011 163 25 250 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=94450 $D=0
M1012 251 26 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=89820 $D=0
M1013 252 26 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=94450 $D=0
M1014 253 249 213 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=89820 $D=0
M1015 254 250 214 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=94450 $D=0
M1016 162 253 699 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=89820 $D=0
M1017 163 254 700 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=94450 $D=0
M1018 255 699 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=89820 $D=0
M1019 256 700 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=94450 $D=0
M1020 253 25 255 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=89820 $D=0
M1021 254 25 256 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=94450 $D=0
M1022 255 251 223 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=89820 $D=0
M1023 256 252 224 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=94450 $D=0
M1024 227 257 255 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=89820 $D=0
M1025 228 258 256 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=94450 $D=0
M1026 257 27 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=89820 $D=0
M1027 258 27 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=94450 $D=0
M1028 162 28 259 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=89820 $D=0
M1029 163 28 260 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=94450 $D=0
M1030 261 29 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=89820 $D=0
M1031 262 29 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=94450 $D=0
M1032 263 259 213 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=89820 $D=0
M1033 264 260 214 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=94450 $D=0
M1034 162 263 701 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=89820 $D=0
M1035 163 264 702 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=94450 $D=0
M1036 265 701 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=89820 $D=0
M1037 266 702 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=94450 $D=0
M1038 263 28 265 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=89820 $D=0
M1039 264 28 266 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=94450 $D=0
M1040 265 261 223 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=89820 $D=0
M1041 266 262 224 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=94450 $D=0
M1042 227 267 265 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=89820 $D=0
M1043 228 268 266 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=94450 $D=0
M1044 267 30 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=89820 $D=0
M1045 268 30 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=94450 $D=0
M1046 162 31 269 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=89820 $D=0
M1047 163 31 270 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=94450 $D=0
M1048 271 32 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=89820 $D=0
M1049 272 32 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=94450 $D=0
M1050 273 269 213 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=89820 $D=0
M1051 274 270 214 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=94450 $D=0
M1052 162 273 703 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=89820 $D=0
M1053 163 274 704 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=94450 $D=0
M1054 275 703 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=89820 $D=0
M1055 276 704 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=94450 $D=0
M1056 273 31 275 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=89820 $D=0
M1057 274 31 276 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=94450 $D=0
M1058 275 271 223 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=89820 $D=0
M1059 276 272 224 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=94450 $D=0
M1060 227 277 275 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=89820 $D=0
M1061 228 278 276 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=94450 $D=0
M1062 277 33 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=89820 $D=0
M1063 278 33 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=94450 $D=0
M1064 162 34 279 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=89820 $D=0
M1065 163 34 280 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=94450 $D=0
M1066 281 35 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=89820 $D=0
M1067 282 35 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=94450 $D=0
M1068 283 279 213 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=89820 $D=0
M1069 284 280 214 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=94450 $D=0
M1070 162 283 705 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=89820 $D=0
M1071 163 284 706 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=94450 $D=0
M1072 285 705 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=89820 $D=0
M1073 286 706 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=94450 $D=0
M1074 283 34 285 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=89820 $D=0
M1075 284 34 286 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=94450 $D=0
M1076 285 281 223 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=89820 $D=0
M1077 286 282 224 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=94450 $D=0
M1078 227 287 285 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=89820 $D=0
M1079 228 288 286 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=94450 $D=0
M1080 287 36 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=89820 $D=0
M1081 288 36 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=94450 $D=0
M1082 162 37 289 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=89820 $D=0
M1083 163 37 290 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=94450 $D=0
M1084 291 38 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=89820 $D=0
M1085 292 38 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=94450 $D=0
M1086 293 289 213 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=89820 $D=0
M1087 294 290 214 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=94450 $D=0
M1088 162 293 707 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=89820 $D=0
M1089 163 294 708 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=94450 $D=0
M1090 295 707 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=89820 $D=0
M1091 296 708 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=94450 $D=0
M1092 293 37 295 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=89820 $D=0
M1093 294 37 296 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=94450 $D=0
M1094 295 291 223 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=89820 $D=0
M1095 296 292 224 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=94450 $D=0
M1096 227 297 295 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=89820 $D=0
M1097 228 298 296 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=94450 $D=0
M1098 297 39 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=89820 $D=0
M1099 298 39 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=94450 $D=0
M1100 162 40 299 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=89820 $D=0
M1101 163 40 300 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=94450 $D=0
M1102 301 41 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=89820 $D=0
M1103 302 41 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=94450 $D=0
M1104 303 299 213 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=89820 $D=0
M1105 304 300 214 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=94450 $D=0
M1106 162 303 709 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=89820 $D=0
M1107 163 304 710 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=94450 $D=0
M1108 305 709 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=89820 $D=0
M1109 306 710 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=94450 $D=0
M1110 303 40 305 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=89820 $D=0
M1111 304 40 306 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=94450 $D=0
M1112 305 301 223 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=89820 $D=0
M1113 306 302 224 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=94450 $D=0
M1114 227 307 305 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=89820 $D=0
M1115 228 308 306 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=94450 $D=0
M1116 307 42 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=89820 $D=0
M1117 308 42 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=94450 $D=0
M1118 162 43 309 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=89820 $D=0
M1119 163 43 310 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=94450 $D=0
M1120 311 44 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=89820 $D=0
M1121 312 44 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=94450 $D=0
M1122 313 309 213 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=89820 $D=0
M1123 314 310 214 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=94450 $D=0
M1124 162 313 711 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=89820 $D=0
M1125 163 314 712 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=94450 $D=0
M1126 315 711 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=89820 $D=0
M1127 316 712 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=94450 $D=0
M1128 313 43 315 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=89820 $D=0
M1129 314 43 316 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=94450 $D=0
M1130 315 311 223 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=89820 $D=0
M1131 316 312 224 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=94450 $D=0
M1132 227 317 315 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=89820 $D=0
M1133 228 318 316 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=94450 $D=0
M1134 317 45 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=89820 $D=0
M1135 318 45 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=94450 $D=0
M1136 162 46 319 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=89820 $D=0
M1137 163 46 320 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=94450 $D=0
M1138 321 47 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=89820 $D=0
M1139 322 47 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=94450 $D=0
M1140 323 319 213 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=89820 $D=0
M1141 324 320 214 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=94450 $D=0
M1142 162 323 713 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=89820 $D=0
M1143 163 324 714 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=94450 $D=0
M1144 325 713 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=89820 $D=0
M1145 326 714 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=94450 $D=0
M1146 323 46 325 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=89820 $D=0
M1147 324 46 326 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=94450 $D=0
M1148 325 321 223 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=89820 $D=0
M1149 326 322 224 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=94450 $D=0
M1150 227 327 325 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=89820 $D=0
M1151 228 328 326 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=94450 $D=0
M1152 327 48 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=89820 $D=0
M1153 328 48 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=94450 $D=0
M1154 162 49 329 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=89820 $D=0
M1155 163 49 330 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=94450 $D=0
M1156 331 50 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=89820 $D=0
M1157 332 50 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=94450 $D=0
M1158 333 329 213 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=89820 $D=0
M1159 334 330 214 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=94450 $D=0
M1160 162 333 715 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=89820 $D=0
M1161 163 334 716 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=94450 $D=0
M1162 335 715 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=89820 $D=0
M1163 336 716 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=94450 $D=0
M1164 333 49 335 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=89820 $D=0
M1165 334 49 336 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=94450 $D=0
M1166 335 331 223 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=89820 $D=0
M1167 336 332 224 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=94450 $D=0
M1168 227 337 335 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=89820 $D=0
M1169 228 338 336 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=94450 $D=0
M1170 337 51 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=89820 $D=0
M1171 338 51 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=94450 $D=0
M1172 162 52 339 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=89820 $D=0
M1173 163 52 340 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=94450 $D=0
M1174 341 53 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=89820 $D=0
M1175 342 53 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=94450 $D=0
M1176 343 339 213 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=89820 $D=0
M1177 344 340 214 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=94450 $D=0
M1178 162 343 717 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=89820 $D=0
M1179 163 344 718 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=94450 $D=0
M1180 345 717 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=89820 $D=0
M1181 346 718 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=94450 $D=0
M1182 343 52 345 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=89820 $D=0
M1183 344 52 346 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=94450 $D=0
M1184 345 341 223 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=89820 $D=0
M1185 346 342 224 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=94450 $D=0
M1186 227 347 345 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=89820 $D=0
M1187 228 348 346 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=94450 $D=0
M1188 347 54 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=89820 $D=0
M1189 348 54 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=94450 $D=0
M1190 162 55 349 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=89820 $D=0
M1191 163 55 350 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=94450 $D=0
M1192 351 56 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=89820 $D=0
M1193 352 56 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=94450 $D=0
M1194 353 349 213 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=89820 $D=0
M1195 354 350 214 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=94450 $D=0
M1196 162 353 719 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=89820 $D=0
M1197 163 354 720 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=94450 $D=0
M1198 355 719 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=89820 $D=0
M1199 356 720 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=94450 $D=0
M1200 353 55 355 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=89820 $D=0
M1201 354 55 356 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=94450 $D=0
M1202 355 351 223 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=89820 $D=0
M1203 356 352 224 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=94450 $D=0
M1204 227 357 355 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=89820 $D=0
M1205 228 358 356 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=94450 $D=0
M1206 357 57 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=89820 $D=0
M1207 358 57 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=94450 $D=0
M1208 162 58 359 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=89820 $D=0
M1209 163 58 360 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=94450 $D=0
M1210 361 59 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=89820 $D=0
M1211 362 59 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=94450 $D=0
M1212 363 359 213 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=89820 $D=0
M1213 364 360 214 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=94450 $D=0
M1214 162 363 721 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=89820 $D=0
M1215 163 364 722 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=94450 $D=0
M1216 365 721 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=89820 $D=0
M1217 366 722 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=94450 $D=0
M1218 363 58 365 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=89820 $D=0
M1219 364 58 366 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=94450 $D=0
M1220 365 361 223 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=89820 $D=0
M1221 366 362 224 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=94450 $D=0
M1222 227 367 365 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=89820 $D=0
M1223 228 368 366 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=94450 $D=0
M1224 367 60 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=89820 $D=0
M1225 368 60 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=94450 $D=0
M1226 162 61 369 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=89820 $D=0
M1227 163 61 370 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=94450 $D=0
M1228 371 62 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=89820 $D=0
M1229 372 62 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=94450 $D=0
M1230 373 369 213 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=89820 $D=0
M1231 374 370 214 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=94450 $D=0
M1232 162 373 723 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=89820 $D=0
M1233 163 374 724 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=94450 $D=0
M1234 375 723 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=89820 $D=0
M1235 376 724 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=94450 $D=0
M1236 373 61 375 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=89820 $D=0
M1237 374 61 376 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=94450 $D=0
M1238 375 371 223 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=89820 $D=0
M1239 376 372 224 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=94450 $D=0
M1240 227 377 375 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=89820 $D=0
M1241 228 378 376 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=94450 $D=0
M1242 377 63 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=89820 $D=0
M1243 378 63 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=94450 $D=0
M1244 162 64 379 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=89820 $D=0
M1245 163 64 380 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=94450 $D=0
M1246 381 65 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=89820 $D=0
M1247 382 65 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=94450 $D=0
M1248 383 379 213 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=89820 $D=0
M1249 384 380 214 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=94450 $D=0
M1250 162 383 725 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=89820 $D=0
M1251 163 384 726 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=94450 $D=0
M1252 385 725 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=89820 $D=0
M1253 386 726 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=94450 $D=0
M1254 383 64 385 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=89820 $D=0
M1255 384 64 386 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=94450 $D=0
M1256 385 381 223 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=89820 $D=0
M1257 386 382 224 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=94450 $D=0
M1258 227 387 385 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=89820 $D=0
M1259 228 388 386 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=94450 $D=0
M1260 387 66 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=89820 $D=0
M1261 388 66 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=94450 $D=0
M1262 162 67 389 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=89820 $D=0
M1263 163 67 390 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=94450 $D=0
M1264 391 68 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=89820 $D=0
M1265 392 68 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=94450 $D=0
M1266 393 389 213 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=89820 $D=0
M1267 394 390 214 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=94450 $D=0
M1268 162 393 727 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=89820 $D=0
M1269 163 394 728 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=94450 $D=0
M1270 395 727 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=89820 $D=0
M1271 396 728 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=94450 $D=0
M1272 393 67 395 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=89820 $D=0
M1273 394 67 396 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=94450 $D=0
M1274 395 391 223 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=89820 $D=0
M1275 396 392 224 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=94450 $D=0
M1276 227 397 395 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=89820 $D=0
M1277 228 398 396 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=94450 $D=0
M1278 397 69 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=89820 $D=0
M1279 398 69 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=94450 $D=0
M1280 162 70 399 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=89820 $D=0
M1281 163 70 400 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=94450 $D=0
M1282 401 71 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=89820 $D=0
M1283 402 71 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=94450 $D=0
M1284 403 399 213 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=89820 $D=0
M1285 404 400 214 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=94450 $D=0
M1286 162 403 729 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=89820 $D=0
M1287 163 404 730 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=94450 $D=0
M1288 405 729 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=89820 $D=0
M1289 406 730 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=94450 $D=0
M1290 403 70 405 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=89820 $D=0
M1291 404 70 406 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=94450 $D=0
M1292 405 401 223 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=89820 $D=0
M1293 406 402 224 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=94450 $D=0
M1294 227 407 405 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=89820 $D=0
M1295 228 408 406 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=94450 $D=0
M1296 407 72 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=89820 $D=0
M1297 408 72 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=94450 $D=0
M1298 162 73 409 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=89820 $D=0
M1299 163 73 410 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=94450 $D=0
M1300 411 74 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=89820 $D=0
M1301 412 74 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=94450 $D=0
M1302 413 409 213 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=89820 $D=0
M1303 414 410 214 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=94450 $D=0
M1304 162 413 731 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=89820 $D=0
M1305 163 414 732 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=94450 $D=0
M1306 415 731 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=89820 $D=0
M1307 416 732 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=94450 $D=0
M1308 413 73 415 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=89820 $D=0
M1309 414 73 416 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=94450 $D=0
M1310 415 411 223 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=89820 $D=0
M1311 416 412 224 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=94450 $D=0
M1312 227 417 415 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=89820 $D=0
M1313 228 418 416 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=94450 $D=0
M1314 417 75 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=89820 $D=0
M1315 418 75 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=94450 $D=0
M1316 162 76 419 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=89820 $D=0
M1317 163 76 420 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=94450 $D=0
M1318 421 77 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=89820 $D=0
M1319 422 77 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=94450 $D=0
M1320 423 419 213 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=89820 $D=0
M1321 424 420 214 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=94450 $D=0
M1322 162 423 733 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=89820 $D=0
M1323 163 424 734 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=94450 $D=0
M1324 425 733 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=89820 $D=0
M1325 426 734 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=94450 $D=0
M1326 423 76 425 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=89820 $D=0
M1327 424 76 426 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=94450 $D=0
M1328 425 421 223 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=89820 $D=0
M1329 426 422 224 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=94450 $D=0
M1330 227 427 425 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=89820 $D=0
M1331 228 428 426 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=94450 $D=0
M1332 427 78 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=89820 $D=0
M1333 428 78 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=94450 $D=0
M1334 162 79 429 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=89820 $D=0
M1335 163 79 430 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=94450 $D=0
M1336 431 80 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=89820 $D=0
M1337 432 80 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=94450 $D=0
M1338 433 429 213 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=89820 $D=0
M1339 434 430 214 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=94450 $D=0
M1340 162 433 735 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=89820 $D=0
M1341 163 434 736 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=94450 $D=0
M1342 435 735 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=89820 $D=0
M1343 436 736 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=94450 $D=0
M1344 433 79 435 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=89820 $D=0
M1345 434 79 436 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=94450 $D=0
M1346 435 431 223 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=89820 $D=0
M1347 436 432 224 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=94450 $D=0
M1348 227 437 435 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=89820 $D=0
M1349 228 438 436 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=94450 $D=0
M1350 437 81 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=89820 $D=0
M1351 438 81 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=94450 $D=0
M1352 162 82 439 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=89820 $D=0
M1353 163 82 440 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=94450 $D=0
M1354 441 83 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=89820 $D=0
M1355 442 83 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=94450 $D=0
M1356 443 439 213 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=89820 $D=0
M1357 444 440 214 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=94450 $D=0
M1358 162 443 737 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=89820 $D=0
M1359 163 444 738 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=94450 $D=0
M1360 445 737 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=89820 $D=0
M1361 446 738 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=94450 $D=0
M1362 443 82 445 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=89820 $D=0
M1363 444 82 446 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=94450 $D=0
M1364 445 441 223 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=89820 $D=0
M1365 446 442 224 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=94450 $D=0
M1366 227 447 445 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=89820 $D=0
M1367 228 448 446 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=94450 $D=0
M1368 447 84 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=89820 $D=0
M1369 448 84 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=94450 $D=0
M1370 162 85 449 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=89820 $D=0
M1371 163 85 450 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=94450 $D=0
M1372 451 86 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=89820 $D=0
M1373 452 86 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=94450 $D=0
M1374 453 449 213 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=89820 $D=0
M1375 454 450 214 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=94450 $D=0
M1376 162 453 739 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=89820 $D=0
M1377 163 454 740 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=94450 $D=0
M1378 455 739 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=89820 $D=0
M1379 456 740 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=94450 $D=0
M1380 453 85 455 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=89820 $D=0
M1381 454 85 456 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=94450 $D=0
M1382 455 451 223 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=89820 $D=0
M1383 456 452 224 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=94450 $D=0
M1384 227 457 455 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=89820 $D=0
M1385 228 458 456 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=94450 $D=0
M1386 457 87 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=89820 $D=0
M1387 458 87 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=94450 $D=0
M1388 162 88 459 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=89820 $D=0
M1389 163 88 460 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=94450 $D=0
M1390 461 89 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=89820 $D=0
M1391 462 89 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=94450 $D=0
M1392 463 459 213 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=89820 $D=0
M1393 464 460 214 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=94450 $D=0
M1394 162 463 741 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=89820 $D=0
M1395 163 464 742 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=94450 $D=0
M1396 465 741 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=89820 $D=0
M1397 466 742 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=94450 $D=0
M1398 463 88 465 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=89820 $D=0
M1399 464 88 466 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=94450 $D=0
M1400 465 461 223 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=89820 $D=0
M1401 466 462 224 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=94450 $D=0
M1402 227 467 465 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=89820 $D=0
M1403 228 468 466 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=94450 $D=0
M1404 467 90 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=89820 $D=0
M1405 468 90 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=94450 $D=0
M1406 162 91 469 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=89820 $D=0
M1407 163 91 470 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=94450 $D=0
M1408 471 92 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=89820 $D=0
M1409 472 92 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=94450 $D=0
M1410 473 469 213 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=89820 $D=0
M1411 474 470 214 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=94450 $D=0
M1412 162 473 743 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=89820 $D=0
M1413 163 474 744 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=94450 $D=0
M1414 475 743 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=89820 $D=0
M1415 476 744 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=94450 $D=0
M1416 473 91 475 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=89820 $D=0
M1417 474 91 476 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=94450 $D=0
M1418 475 471 223 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=89820 $D=0
M1419 476 472 224 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=94450 $D=0
M1420 227 477 475 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=89820 $D=0
M1421 228 478 476 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=94450 $D=0
M1422 477 93 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=89820 $D=0
M1423 478 93 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=94450 $D=0
M1424 162 94 479 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=89820 $D=0
M1425 163 94 480 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=94450 $D=0
M1426 481 95 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=89820 $D=0
M1427 482 95 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=94450 $D=0
M1428 483 479 213 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=89820 $D=0
M1429 484 480 214 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=94450 $D=0
M1430 162 483 745 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=89820 $D=0
M1431 163 484 746 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=94450 $D=0
M1432 485 745 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=89820 $D=0
M1433 486 746 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=94450 $D=0
M1434 483 94 485 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=89820 $D=0
M1435 484 94 486 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=94450 $D=0
M1436 485 481 223 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=89820 $D=0
M1437 486 482 224 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=94450 $D=0
M1438 227 487 485 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=89820 $D=0
M1439 228 488 486 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=94450 $D=0
M1440 487 96 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=89820 $D=0
M1441 488 96 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=94450 $D=0
M1442 162 97 489 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=89820 $D=0
M1443 163 97 490 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=94450 $D=0
M1444 491 98 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=89820 $D=0
M1445 492 98 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=94450 $D=0
M1446 493 489 213 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=89820 $D=0
M1447 494 490 214 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=94450 $D=0
M1448 162 493 747 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=89820 $D=0
M1449 163 494 748 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=94450 $D=0
M1450 495 747 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=89820 $D=0
M1451 496 748 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=94450 $D=0
M1452 493 97 495 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=89820 $D=0
M1453 494 97 496 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=94450 $D=0
M1454 495 491 223 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=89820 $D=0
M1455 496 492 224 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=94450 $D=0
M1456 227 497 495 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=89820 $D=0
M1457 228 498 496 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=94450 $D=0
M1458 497 99 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=89820 $D=0
M1459 498 99 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=94450 $D=0
M1460 162 100 499 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=89820 $D=0
M1461 163 100 500 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=94450 $D=0
M1462 501 101 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=89820 $D=0
M1463 502 101 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=94450 $D=0
M1464 503 499 213 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=89820 $D=0
M1465 504 500 214 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=94450 $D=0
M1466 162 503 749 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=89820 $D=0
M1467 163 504 750 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=94450 $D=0
M1468 505 749 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=89820 $D=0
M1469 506 750 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=94450 $D=0
M1470 503 100 505 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=89820 $D=0
M1471 504 100 506 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=94450 $D=0
M1472 505 501 223 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=89820 $D=0
M1473 506 502 224 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=94450 $D=0
M1474 227 507 505 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=89820 $D=0
M1475 228 508 506 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=94450 $D=0
M1476 507 102 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=89820 $D=0
M1477 508 102 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=94450 $D=0
M1478 162 103 509 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=89820 $D=0
M1479 163 103 510 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=94450 $D=0
M1480 511 104 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=89820 $D=0
M1481 512 104 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=94450 $D=0
M1482 513 509 213 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=89820 $D=0
M1483 514 510 214 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=94450 $D=0
M1484 162 513 751 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=89820 $D=0
M1485 163 514 752 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=94450 $D=0
M1486 515 751 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=89820 $D=0
M1487 516 752 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=94450 $D=0
M1488 513 103 515 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=89820 $D=0
M1489 514 103 516 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=94450 $D=0
M1490 515 511 223 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=89820 $D=0
M1491 516 512 224 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=94450 $D=0
M1492 227 517 515 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=89820 $D=0
M1493 228 518 516 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=94450 $D=0
M1494 517 105 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=89820 $D=0
M1495 518 105 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=94450 $D=0
M1496 162 106 519 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=89820 $D=0
M1497 163 106 520 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=94450 $D=0
M1498 521 107 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=89820 $D=0
M1499 522 107 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=94450 $D=0
M1500 523 519 213 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=89820 $D=0
M1501 524 520 214 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=94450 $D=0
M1502 162 523 753 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=89820 $D=0
M1503 163 524 754 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=94450 $D=0
M1504 525 753 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=89820 $D=0
M1505 526 754 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=94450 $D=0
M1506 523 106 525 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=89820 $D=0
M1507 524 106 526 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=94450 $D=0
M1508 525 521 223 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=89820 $D=0
M1509 526 522 224 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=94450 $D=0
M1510 227 527 525 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=89820 $D=0
M1511 228 528 526 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=94450 $D=0
M1512 527 108 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=89820 $D=0
M1513 528 108 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=94450 $D=0
M1514 162 109 529 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=89820 $D=0
M1515 163 109 530 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=94450 $D=0
M1516 531 110 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=89820 $D=0
M1517 532 110 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=94450 $D=0
M1518 5 531 223 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=89820 $D=0
M1519 6 532 224 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=94450 $D=0
M1520 227 529 5 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=89820 $D=0
M1521 228 530 6 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=94450 $D=0
M1522 162 535 533 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=89820 $D=0
M1523 163 536 534 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=94450 $D=0
M1524 535 111 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=89820 $D=0
M1525 536 111 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=94450 $D=0
M1526 755 223 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=89820 $D=0
M1527 756 224 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=94450 $D=0
M1528 537 535 755 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=89820 $D=0
M1529 538 536 756 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=94450 $D=0
M1530 162 537 539 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=89820 $D=0
M1531 163 538 540 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=94450 $D=0
M1532 757 539 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=89820 $D=0
M1533 758 540 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=94450 $D=0
M1534 537 533 757 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=89820 $D=0
M1535 538 534 758 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=94450 $D=0
M1536 162 543 541 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=89820 $D=0
M1537 163 544 542 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=94450 $D=0
M1538 543 111 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=89820 $D=0
M1539 544 111 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=94450 $D=0
M1540 759 227 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=89820 $D=0
M1541 760 228 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=94450 $D=0
M1542 545 543 759 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=89820 $D=0
M1543 546 544 760 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=94450 $D=0
M1544 162 545 112 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=89820 $D=0
M1545 163 546 113 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=94450 $D=0
M1546 761 112 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=89820 $D=0
M1547 762 113 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=94450 $D=0
M1548 545 541 761 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=89820 $D=0
M1549 546 542 762 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=94450 $D=0
M1550 547 114 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=89820 $D=0
M1551 548 114 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=94450 $D=0
M1552 549 114 539 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=89820 $D=0
M1553 550 114 540 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=94450 $D=0
M1554 115 547 549 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=89820 $D=0
M1555 116 548 550 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=94450 $D=0
M1556 551 117 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=89820 $D=0
M1557 552 117 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=94450 $D=0
M1558 553 117 112 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=89820 $D=0
M1559 554 117 113 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=94450 $D=0
M1560 763 551 553 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=89820 $D=0
M1561 764 552 554 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=94450 $D=0
M1562 162 112 763 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=89820 $D=0
M1563 163 113 764 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=94450 $D=0
M1564 555 118 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=89820 $D=0
M1565 556 118 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=94450 $D=0
M1566 557 118 553 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=89820 $D=0
M1567 558 118 554 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=94450 $D=0
M1568 10 555 557 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=89820 $D=0
M1569 11 556 558 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=94450 $D=0
M1570 560 559 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=89820 $D=0
M1571 561 119 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=94450 $D=0
M1572 162 564 562 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=89820 $D=0
M1573 163 565 563 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=94450 $D=0
M1574 566 549 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=89820 $D=0
M1575 567 550 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=94450 $D=0
M1576 564 549 559 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=89820 $D=0
M1577 565 550 119 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=94450 $D=0
M1578 560 566 564 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=89820 $D=0
M1579 561 567 565 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=94450 $D=0
M1580 568 562 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=89820 $D=0
M1581 569 563 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=94450 $D=0
M1582 570 562 557 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=89820 $D=0
M1583 559 563 558 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=94450 $D=0
M1584 549 568 570 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=89820 $D=0
M1585 550 569 559 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=94450 $D=0
M1586 571 570 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=89820 $D=0
M1587 572 559 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=94450 $D=0
M1588 573 562 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=89820 $D=0
M1589 574 563 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=94450 $D=0
M1590 575 562 571 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=89820 $D=0
M1591 576 563 572 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=94450 $D=0
M1592 557 573 575 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=89820 $D=0
M1593 558 574 576 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=94450 $D=0
M1594 786 549 162 162 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=89460 $D=0
M1595 787 550 163 163 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=94090 $D=0
M1596 577 557 786 162 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=89460 $D=0
M1597 578 558 787 163 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=94090 $D=0
M1598 579 575 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=89820 $D=0
M1599 580 576 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=94450 $D=0
M1600 581 549 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=89820 $D=0
M1601 582 550 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=94450 $D=0
M1602 162 557 581 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=89820 $D=0
M1603 163 558 582 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=94450 $D=0
M1604 583 549 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=89820 $D=0
M1605 584 550 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=94450 $D=0
M1606 162 557 583 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=89820 $D=0
M1607 163 558 584 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=94450 $D=0
M1608 788 549 162 162 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=89640 $D=0
M1609 789 550 163 163 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=94270 $D=0
M1610 587 557 788 162 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=89640 $D=0
M1611 588 558 789 163 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=94270 $D=0
M1612 162 583 587 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=89820 $D=0
M1613 163 584 588 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=94450 $D=0
M1614 589 121 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=89820 $D=0
M1615 590 121 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=94450 $D=0
M1616 591 121 577 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=89820 $D=0
M1617 592 121 578 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=94450 $D=0
M1618 581 589 591 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=89820 $D=0
M1619 582 590 592 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=94450 $D=0
M1620 593 121 579 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=89820 $D=0
M1621 594 121 580 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=94450 $D=0
M1622 587 589 593 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=89820 $D=0
M1623 588 590 594 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=94450 $D=0
M1624 595 122 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=89820 $D=0
M1625 596 122 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=94450 $D=0
M1626 597 122 593 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=89820 $D=0
M1627 598 122 594 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=94450 $D=0
M1628 591 595 597 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=89820 $D=0
M1629 592 596 598 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=94450 $D=0
M1630 12 597 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=89820 $D=0
M1631 13 598 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=94450 $D=0
M1632 599 123 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=89820 $D=0
M1633 600 123 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=94450 $D=0
M1634 601 123 124 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=89820 $D=0
M1635 602 123 125 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=94450 $D=0
M1636 126 599 601 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=89820 $D=0
M1637 127 600 602 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=94450 $D=0
M1638 603 123 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=89820 $D=0
M1639 604 123 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=94450 $D=0
M1640 609 123 128 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=89820 $D=0
M1641 610 123 130 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=94450 $D=0
M1642 131 603 609 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=89820 $D=0
M1643 129 604 610 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=94450 $D=0
M1644 611 123 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=89820 $D=0
M1645 612 123 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=94450 $D=0
M1646 613 123 132 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=89820 $D=0
M1647 614 123 133 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=94450 $D=0
M1648 134 611 613 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=89820 $D=0
M1649 135 612 614 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=94450 $D=0
M1650 615 123 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=89820 $D=0
M1651 616 123 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=94450 $D=0
M1652 617 123 136 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=89820 $D=0
M1653 618 123 137 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=94450 $D=0
M1654 138 615 617 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=89820 $D=0
M1655 139 616 618 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=94450 $D=0
M1656 619 123 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=89820 $D=0
M1657 620 123 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=94450 $D=0
M1658 621 123 5 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=89820 $D=0
M1659 622 123 6 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=94450 $D=0
M1660 140 619 621 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=89820 $D=0
M1661 141 620 622 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=94450 $D=0
M1662 162 549 776 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=89820 $D=0
M1663 163 550 777 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=94450 $D=0
M1664 127 776 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=89820 $D=0
M1665 124 777 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=94450 $D=0
M1666 623 142 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=89820 $D=0
M1667 624 142 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=94450 $D=0
M1668 143 142 127 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=89820 $D=0
M1669 144 142 124 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=94450 $D=0
M1670 601 623 143 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=89820 $D=0
M1671 602 624 144 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=94450 $D=0
M1672 625 145 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=89820 $D=0
M1673 626 145 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=94450 $D=0
M1674 120 145 143 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=89820 $D=0
M1675 146 145 144 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=94450 $D=0
M1676 609 625 120 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=89820 $D=0
M1677 610 626 146 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=94450 $D=0
M1678 627 147 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=89820 $D=0
M1679 628 147 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=94450 $D=0
M1680 148 147 120 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=89820 $D=0
M1681 149 147 146 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=94450 $D=0
M1682 613 627 148 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=89820 $D=0
M1683 614 628 149 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=94450 $D=0
M1684 629 150 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=89820 $D=0
M1685 630 150 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=94450 $D=0
M1686 151 150 148 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=89820 $D=0
M1687 152 150 149 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=94450 $D=0
M1688 617 629 151 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=89820 $D=0
M1689 618 630 152 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=94450 $D=0
M1690 631 153 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=89820 $D=0
M1691 632 153 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=94450 $D=0
M1692 199 153 151 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=89820 $D=0
M1693 200 153 152 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=94450 $D=0
M1694 621 631 199 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=89820 $D=0
M1695 622 632 200 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=94450 $D=0
M1696 633 154 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=89820 $D=0
M1697 634 154 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=94450 $D=0
M1698 635 154 112 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=89820 $D=0
M1699 636 154 113 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=94450 $D=0
M1700 10 633 635 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=89820 $D=0
M1701 11 634 636 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=94450 $D=0
M1702 637 539 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=89820 $D=0
M1703 638 540 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=94450 $D=0
M1704 162 635 637 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=89820 $D=0
M1705 163 636 638 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=94450 $D=0
M1706 790 539 162 162 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=89640 $D=0
M1707 791 540 163 163 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=94270 $D=0
M1708 641 635 790 162 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=89640 $D=0
M1709 642 636 791 163 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=94270 $D=0
M1710 162 637 641 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=89820 $D=0
M1711 163 638 642 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=94450 $D=0
M1712 778 643 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=89820 $D=0
M1713 779 644 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=94450 $D=0
M1714 162 641 778 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=89820 $D=0
M1715 163 642 779 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=94450 $D=0
M1716 644 778 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=89820 $D=0
M1717 155 779 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=94450 $D=0
M1718 792 539 162 162 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=89460 $D=0
M1719 793 540 163 163 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=94090 $D=0
M1720 645 647 792 162 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=89460 $D=0
M1721 646 648 793 163 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=94090 $D=0
M1722 647 635 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=89820 $D=0
M1723 648 636 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=94450 $D=0
M1724 649 645 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=89820 $D=0
M1725 650 646 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=94450 $D=0
M1726 162 643 649 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=89820 $D=0
M1727 163 644 650 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=94450 $D=0
M1728 652 156 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=89820 $D=0
M1729 653 651 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=94450 $D=0
M1730 651 649 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=89820 $D=0
M1731 157 650 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=94450 $D=0
M1732 162 652 651 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=89820 $D=0
M1733 163 653 157 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=94450 $D=0
M1734 655 654 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=89820 $D=0
M1735 656 158 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=94450 $D=0
M1736 162 659 657 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=89820 $D=0
M1737 163 660 658 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=94450 $D=0
M1738 661 115 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=89820 $D=0
M1739 662 116 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=94450 $D=0
M1740 659 115 654 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=89820 $D=0
M1741 660 116 158 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=94450 $D=0
M1742 655 661 659 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=89820 $D=0
M1743 656 662 660 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=94450 $D=0
M1744 663 657 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=89820 $D=0
M1745 664 658 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=94450 $D=0
M1746 159 657 5 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=89820 $D=0
M1747 654 658 6 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=94450 $D=0
M1748 115 663 159 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=89820 $D=0
M1749 116 664 654 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=94450 $D=0
M1750 665 159 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=89820 $D=0
M1751 666 654 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=94450 $D=0
M1752 667 657 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=89820 $D=0
M1753 668 658 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=94450 $D=0
M1754 201 657 665 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=89820 $D=0
M1755 202 658 666 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=94450 $D=0
M1756 5 667 201 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=89820 $D=0
M1757 6 668 202 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=94450 $D=0
M1758 669 160 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=89820 $D=0
M1759 670 160 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=94450 $D=0
M1760 671 160 201 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=89820 $D=0
M1761 672 160 202 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=94450 $D=0
M1762 12 669 671 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=89820 $D=0
M1763 13 670 672 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=94450 $D=0
M1764 673 161 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=89820 $D=0
M1765 674 161 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=94450 $D=0
M1766 161 161 671 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=89820 $D=0
M1767 161 161 672 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=94450 $D=0
M1768 5 673 161 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=89820 $D=0
M1769 6 674 161 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=94450 $D=0
M1770 675 111 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=89820 $D=0
M1771 676 111 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=94450 $D=0
M1772 162 675 677 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=89820 $D=0
M1773 163 676 678 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=94450 $D=0
M1774 679 111 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=89820 $D=0
M1775 680 111 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=94450 $D=0
M1776 681 677 161 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=89820 $D=0
M1777 682 678 161 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=94450 $D=0
M1778 162 681 780 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=89820 $D=0
M1779 163 682 781 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=94450 $D=0
M1780 683 780 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=89820 $D=0
M1781 684 781 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=94450 $D=0
M1782 681 675 683 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=89820 $D=0
M1783 682 676 684 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=94450 $D=0
M1784 685 679 683 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=89820 $D=0
M1785 686 680 684 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=94450 $D=0
M1786 162 689 687 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=89820 $D=0
M1787 163 690 688 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=94450 $D=0
M1788 689 111 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=89820 $D=0
M1789 690 111 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=94450 $D=0
M1790 782 685 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=89820 $D=0
M1791 783 686 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=94450 $D=0
M1792 691 689 782 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=89820 $D=0
M1793 692 690 783 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=94450 $D=0
M1794 162 691 115 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=89820 $D=0
M1795 163 692 116 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=94450 $D=0
M1796 784 115 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=89820 $D=0
M1797 785 116 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=94450 $D=0
M1798 691 687 784 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=89820 $D=0
M1799 692 688 785 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=94450 $D=0
.ENDS
***************************************
.SUBCKT ICV_30 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164
** N=801 EP=164 IP=1514 FDC=1800
M0 174 1 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=79310 $D=1
M1 175 1 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=83940 $D=1
M2 176 174 2 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=79310 $D=1
M3 177 175 3 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=83940 $D=1
M4 5 1 176 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=79310 $D=1
M5 6 1 177 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=83940 $D=1
M6 178 174 4 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=79310 $D=1
M7 179 175 4 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=83940 $D=1
M8 2 1 178 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=79310 $D=1
M9 3 1 179 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=83940 $D=1
M10 180 174 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=79310 $D=1
M11 181 175 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=83940 $D=1
M12 2 1 180 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=79310 $D=1
M13 3 1 181 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=83940 $D=1
M14 184 182 180 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=79310 $D=1
M15 185 183 181 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=83940 $D=1
M16 182 7 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=79310 $D=1
M17 183 7 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=83940 $D=1
M18 186 182 178 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=79310 $D=1
M19 187 183 179 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=83940 $D=1
M20 176 7 186 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=79310 $D=1
M21 177 7 187 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=83940 $D=1
M22 188 8 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=79310 $D=1
M23 189 8 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=83940 $D=1
M24 190 188 186 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=79310 $D=1
M25 191 189 187 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=83940 $D=1
M26 184 8 190 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=79310 $D=1
M27 185 8 191 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=83940 $D=1
M28 192 9 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=79310 $D=1
M29 193 9 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=83940 $D=1
M30 194 192 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=79310 $D=1
M31 195 193 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=83940 $D=1
M32 10 9 194 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=79310 $D=1
M33 11 9 195 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=83940 $D=1
M34 196 192 12 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=79310 $D=1
M35 197 193 13 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=83940 $D=1
M36 198 9 196 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=79310 $D=1
M37 199 9 197 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=83940 $D=1
M38 202 192 200 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=79310 $D=1
M39 203 193 201 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=83940 $D=1
M40 190 9 202 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=79310 $D=1
M41 191 9 203 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=83940 $D=1
M42 206 204 202 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=79310 $D=1
M43 207 205 203 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=83940 $D=1
M44 204 14 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=79310 $D=1
M45 205 14 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=83940 $D=1
M46 208 204 196 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=79310 $D=1
M47 209 205 197 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=83940 $D=1
M48 194 14 208 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=79310 $D=1
M49 195 14 209 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=83940 $D=1
M50 210 15 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=79310 $D=1
M51 211 15 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=83940 $D=1
M52 212 210 208 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=79310 $D=1
M53 213 211 209 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=83940 $D=1
M54 206 15 212 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=79310 $D=1
M55 207 15 213 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=83940 $D=1
M56 5 16 214 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=79310 $D=1
M57 6 16 215 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=83940 $D=1
M58 216 17 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=79310 $D=1
M59 217 17 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=83940 $D=1
M60 218 16 212 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=79310 $D=1
M61 219 16 213 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=83940 $D=1
M62 5 218 690 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=79310 $D=1
M63 6 219 691 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=83940 $D=1
M64 220 690 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=79310 $D=1
M65 221 691 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=83940 $D=1
M66 218 214 220 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=79310 $D=1
M67 219 215 221 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=83940 $D=1
M68 220 17 222 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=79310 $D=1
M69 221 17 223 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=83940 $D=1
M70 226 18 220 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=79310 $D=1
M71 227 18 221 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=83940 $D=1
M72 224 18 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=79310 $D=1
M73 225 18 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=83940 $D=1
M74 5 19 228 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=79310 $D=1
M75 6 19 229 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=83940 $D=1
M76 230 20 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=79310 $D=1
M77 231 20 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=83940 $D=1
M78 232 19 212 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=79310 $D=1
M79 233 19 213 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=83940 $D=1
M80 5 232 692 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=79310 $D=1
M81 6 233 693 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=83940 $D=1
M82 234 692 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=79310 $D=1
M83 235 693 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=83940 $D=1
M84 232 228 234 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=79310 $D=1
M85 233 229 235 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=83940 $D=1
M86 234 20 222 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=79310 $D=1
M87 235 20 223 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=83940 $D=1
M88 226 21 234 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=79310 $D=1
M89 227 21 235 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=83940 $D=1
M90 236 21 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=79310 $D=1
M91 237 21 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=83940 $D=1
M92 5 22 238 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=79310 $D=1
M93 6 22 239 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=83940 $D=1
M94 240 23 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=79310 $D=1
M95 241 23 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=83940 $D=1
M96 242 22 212 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=79310 $D=1
M97 243 22 213 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=83940 $D=1
M98 5 242 694 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=79310 $D=1
M99 6 243 695 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=83940 $D=1
M100 244 694 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=79310 $D=1
M101 245 695 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=83940 $D=1
M102 242 238 244 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=79310 $D=1
M103 243 239 245 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=83940 $D=1
M104 244 23 222 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=79310 $D=1
M105 245 23 223 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=83940 $D=1
M106 226 24 244 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=79310 $D=1
M107 227 24 245 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=83940 $D=1
M108 246 24 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=79310 $D=1
M109 247 24 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=83940 $D=1
M110 5 25 248 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=79310 $D=1
M111 6 25 249 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=83940 $D=1
M112 250 26 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=79310 $D=1
M113 251 26 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=83940 $D=1
M114 252 25 212 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=79310 $D=1
M115 253 25 213 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=83940 $D=1
M116 5 252 696 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=79310 $D=1
M117 6 253 697 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=83940 $D=1
M118 254 696 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=79310 $D=1
M119 255 697 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=83940 $D=1
M120 252 248 254 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=79310 $D=1
M121 253 249 255 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=83940 $D=1
M122 254 26 222 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=79310 $D=1
M123 255 26 223 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=83940 $D=1
M124 226 27 254 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=79310 $D=1
M125 227 27 255 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=83940 $D=1
M126 256 27 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=79310 $D=1
M127 257 27 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=83940 $D=1
M128 5 28 258 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=79310 $D=1
M129 6 28 259 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=83940 $D=1
M130 260 29 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=79310 $D=1
M131 261 29 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=83940 $D=1
M132 262 28 212 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=79310 $D=1
M133 263 28 213 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=83940 $D=1
M134 5 262 698 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=79310 $D=1
M135 6 263 699 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=83940 $D=1
M136 264 698 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=79310 $D=1
M137 265 699 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=83940 $D=1
M138 262 258 264 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=79310 $D=1
M139 263 259 265 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=83940 $D=1
M140 264 29 222 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=79310 $D=1
M141 265 29 223 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=83940 $D=1
M142 226 30 264 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=79310 $D=1
M143 227 30 265 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=83940 $D=1
M144 266 30 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=79310 $D=1
M145 267 30 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=83940 $D=1
M146 5 31 268 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=79310 $D=1
M147 6 31 269 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=83940 $D=1
M148 270 32 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=79310 $D=1
M149 271 32 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=83940 $D=1
M150 272 31 212 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=79310 $D=1
M151 273 31 213 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=83940 $D=1
M152 5 272 700 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=79310 $D=1
M153 6 273 701 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=83940 $D=1
M154 274 700 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=79310 $D=1
M155 275 701 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=83940 $D=1
M156 272 268 274 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=79310 $D=1
M157 273 269 275 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=83940 $D=1
M158 274 32 222 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=79310 $D=1
M159 275 32 223 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=83940 $D=1
M160 226 33 274 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=79310 $D=1
M161 227 33 275 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=83940 $D=1
M162 276 33 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=79310 $D=1
M163 277 33 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=83940 $D=1
M164 5 34 278 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=79310 $D=1
M165 6 34 279 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=83940 $D=1
M166 280 35 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=79310 $D=1
M167 281 35 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=83940 $D=1
M168 282 34 212 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=79310 $D=1
M169 283 34 213 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=83940 $D=1
M170 5 282 702 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=79310 $D=1
M171 6 283 703 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=83940 $D=1
M172 284 702 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=79310 $D=1
M173 285 703 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=83940 $D=1
M174 282 278 284 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=79310 $D=1
M175 283 279 285 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=83940 $D=1
M176 284 35 222 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=79310 $D=1
M177 285 35 223 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=83940 $D=1
M178 226 36 284 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=79310 $D=1
M179 227 36 285 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=83940 $D=1
M180 286 36 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=79310 $D=1
M181 287 36 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=83940 $D=1
M182 5 37 288 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=79310 $D=1
M183 6 37 289 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=83940 $D=1
M184 290 38 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=79310 $D=1
M185 291 38 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=83940 $D=1
M186 292 37 212 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=79310 $D=1
M187 293 37 213 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=83940 $D=1
M188 5 292 704 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=79310 $D=1
M189 6 293 705 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=83940 $D=1
M190 294 704 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=79310 $D=1
M191 295 705 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=83940 $D=1
M192 292 288 294 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=79310 $D=1
M193 293 289 295 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=83940 $D=1
M194 294 38 222 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=79310 $D=1
M195 295 38 223 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=83940 $D=1
M196 226 39 294 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=79310 $D=1
M197 227 39 295 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=83940 $D=1
M198 296 39 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=79310 $D=1
M199 297 39 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=83940 $D=1
M200 5 40 298 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=79310 $D=1
M201 6 40 299 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=83940 $D=1
M202 300 41 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=79310 $D=1
M203 301 41 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=83940 $D=1
M204 302 40 212 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=79310 $D=1
M205 303 40 213 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=83940 $D=1
M206 5 302 706 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=79310 $D=1
M207 6 303 707 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=83940 $D=1
M208 304 706 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=79310 $D=1
M209 305 707 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=83940 $D=1
M210 302 298 304 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=79310 $D=1
M211 303 299 305 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=83940 $D=1
M212 304 41 222 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=79310 $D=1
M213 305 41 223 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=83940 $D=1
M214 226 42 304 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=79310 $D=1
M215 227 42 305 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=83940 $D=1
M216 306 42 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=79310 $D=1
M217 307 42 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=83940 $D=1
M218 5 43 308 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=79310 $D=1
M219 6 43 309 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=83940 $D=1
M220 310 44 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=79310 $D=1
M221 311 44 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=83940 $D=1
M222 312 43 212 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=79310 $D=1
M223 313 43 213 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=83940 $D=1
M224 5 312 708 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=79310 $D=1
M225 6 313 709 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=83940 $D=1
M226 314 708 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=79310 $D=1
M227 315 709 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=83940 $D=1
M228 312 308 314 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=79310 $D=1
M229 313 309 315 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=83940 $D=1
M230 314 44 222 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=79310 $D=1
M231 315 44 223 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=83940 $D=1
M232 226 45 314 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=79310 $D=1
M233 227 45 315 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=83940 $D=1
M234 316 45 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=79310 $D=1
M235 317 45 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=83940 $D=1
M236 5 46 318 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=79310 $D=1
M237 6 46 319 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=83940 $D=1
M238 320 47 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=79310 $D=1
M239 321 47 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=83940 $D=1
M240 322 46 212 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=79310 $D=1
M241 323 46 213 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=83940 $D=1
M242 5 322 710 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=79310 $D=1
M243 6 323 711 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=83940 $D=1
M244 324 710 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=79310 $D=1
M245 325 711 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=83940 $D=1
M246 322 318 324 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=79310 $D=1
M247 323 319 325 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=83940 $D=1
M248 324 47 222 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=79310 $D=1
M249 325 47 223 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=83940 $D=1
M250 226 48 324 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=79310 $D=1
M251 227 48 325 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=83940 $D=1
M252 326 48 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=79310 $D=1
M253 327 48 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=83940 $D=1
M254 5 49 328 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=79310 $D=1
M255 6 49 329 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=83940 $D=1
M256 330 50 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=79310 $D=1
M257 331 50 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=83940 $D=1
M258 332 49 212 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=79310 $D=1
M259 333 49 213 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=83940 $D=1
M260 5 332 712 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=79310 $D=1
M261 6 333 713 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=83940 $D=1
M262 334 712 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=79310 $D=1
M263 335 713 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=83940 $D=1
M264 332 328 334 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=79310 $D=1
M265 333 329 335 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=83940 $D=1
M266 334 50 222 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=79310 $D=1
M267 335 50 223 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=83940 $D=1
M268 226 51 334 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=79310 $D=1
M269 227 51 335 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=83940 $D=1
M270 336 51 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=79310 $D=1
M271 337 51 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=83940 $D=1
M272 5 52 338 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=79310 $D=1
M273 6 52 339 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=83940 $D=1
M274 340 53 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=79310 $D=1
M275 341 53 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=83940 $D=1
M276 342 52 212 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=79310 $D=1
M277 343 52 213 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=83940 $D=1
M278 5 342 714 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=79310 $D=1
M279 6 343 715 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=83940 $D=1
M280 344 714 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=79310 $D=1
M281 345 715 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=83940 $D=1
M282 342 338 344 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=79310 $D=1
M283 343 339 345 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=83940 $D=1
M284 344 53 222 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=79310 $D=1
M285 345 53 223 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=83940 $D=1
M286 226 54 344 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=79310 $D=1
M287 227 54 345 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=83940 $D=1
M288 346 54 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=79310 $D=1
M289 347 54 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=83940 $D=1
M290 5 55 348 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=79310 $D=1
M291 6 55 349 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=83940 $D=1
M292 350 56 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=79310 $D=1
M293 351 56 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=83940 $D=1
M294 352 55 212 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=79310 $D=1
M295 353 55 213 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=83940 $D=1
M296 5 352 716 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=79310 $D=1
M297 6 353 717 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=83940 $D=1
M298 354 716 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=79310 $D=1
M299 355 717 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=83940 $D=1
M300 352 348 354 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=79310 $D=1
M301 353 349 355 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=83940 $D=1
M302 354 56 222 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=79310 $D=1
M303 355 56 223 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=83940 $D=1
M304 226 57 354 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=79310 $D=1
M305 227 57 355 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=83940 $D=1
M306 356 57 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=79310 $D=1
M307 357 57 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=83940 $D=1
M308 5 58 358 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=79310 $D=1
M309 6 58 359 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=83940 $D=1
M310 360 59 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=79310 $D=1
M311 361 59 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=83940 $D=1
M312 362 58 212 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=79310 $D=1
M313 363 58 213 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=83940 $D=1
M314 5 362 718 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=79310 $D=1
M315 6 363 719 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=83940 $D=1
M316 364 718 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=79310 $D=1
M317 365 719 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=83940 $D=1
M318 362 358 364 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=79310 $D=1
M319 363 359 365 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=83940 $D=1
M320 364 59 222 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=79310 $D=1
M321 365 59 223 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=83940 $D=1
M322 226 60 364 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=79310 $D=1
M323 227 60 365 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=83940 $D=1
M324 366 60 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=79310 $D=1
M325 367 60 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=83940 $D=1
M326 5 61 368 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=79310 $D=1
M327 6 61 369 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=83940 $D=1
M328 370 62 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=79310 $D=1
M329 371 62 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=83940 $D=1
M330 372 61 212 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=79310 $D=1
M331 373 61 213 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=83940 $D=1
M332 5 372 720 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=79310 $D=1
M333 6 373 721 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=83940 $D=1
M334 374 720 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=79310 $D=1
M335 375 721 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=83940 $D=1
M336 372 368 374 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=79310 $D=1
M337 373 369 375 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=83940 $D=1
M338 374 62 222 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=79310 $D=1
M339 375 62 223 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=83940 $D=1
M340 226 63 374 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=79310 $D=1
M341 227 63 375 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=83940 $D=1
M342 376 63 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=79310 $D=1
M343 377 63 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=83940 $D=1
M344 5 64 378 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=79310 $D=1
M345 6 64 379 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=83940 $D=1
M346 380 65 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=79310 $D=1
M347 381 65 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=83940 $D=1
M348 382 64 212 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=79310 $D=1
M349 383 64 213 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=83940 $D=1
M350 5 382 722 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=79310 $D=1
M351 6 383 723 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=83940 $D=1
M352 384 722 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=79310 $D=1
M353 385 723 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=83940 $D=1
M354 382 378 384 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=79310 $D=1
M355 383 379 385 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=83940 $D=1
M356 384 65 222 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=79310 $D=1
M357 385 65 223 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=83940 $D=1
M358 226 66 384 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=79310 $D=1
M359 227 66 385 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=83940 $D=1
M360 386 66 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=79310 $D=1
M361 387 66 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=83940 $D=1
M362 5 67 388 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=79310 $D=1
M363 6 67 389 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=83940 $D=1
M364 390 68 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=79310 $D=1
M365 391 68 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=83940 $D=1
M366 392 67 212 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=79310 $D=1
M367 393 67 213 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=83940 $D=1
M368 5 392 724 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=79310 $D=1
M369 6 393 725 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=83940 $D=1
M370 394 724 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=79310 $D=1
M371 395 725 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=83940 $D=1
M372 392 388 394 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=79310 $D=1
M373 393 389 395 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=83940 $D=1
M374 394 68 222 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=79310 $D=1
M375 395 68 223 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=83940 $D=1
M376 226 69 394 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=79310 $D=1
M377 227 69 395 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=83940 $D=1
M378 396 69 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=79310 $D=1
M379 397 69 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=83940 $D=1
M380 5 70 398 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=79310 $D=1
M381 6 70 399 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=83940 $D=1
M382 400 71 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=79310 $D=1
M383 401 71 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=83940 $D=1
M384 402 70 212 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=79310 $D=1
M385 403 70 213 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=83940 $D=1
M386 5 402 726 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=79310 $D=1
M387 6 403 727 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=83940 $D=1
M388 404 726 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=79310 $D=1
M389 405 727 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=83940 $D=1
M390 402 398 404 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=79310 $D=1
M391 403 399 405 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=83940 $D=1
M392 404 71 222 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=79310 $D=1
M393 405 71 223 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=83940 $D=1
M394 226 72 404 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=79310 $D=1
M395 227 72 405 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=83940 $D=1
M396 406 72 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=79310 $D=1
M397 407 72 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=83940 $D=1
M398 5 73 408 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=79310 $D=1
M399 6 73 409 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=83940 $D=1
M400 410 74 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=79310 $D=1
M401 411 74 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=83940 $D=1
M402 412 73 212 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=79310 $D=1
M403 413 73 213 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=83940 $D=1
M404 5 412 728 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=79310 $D=1
M405 6 413 729 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=83940 $D=1
M406 414 728 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=79310 $D=1
M407 415 729 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=83940 $D=1
M408 412 408 414 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=79310 $D=1
M409 413 409 415 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=83940 $D=1
M410 414 74 222 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=79310 $D=1
M411 415 74 223 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=83940 $D=1
M412 226 75 414 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=79310 $D=1
M413 227 75 415 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=83940 $D=1
M414 416 75 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=79310 $D=1
M415 417 75 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=83940 $D=1
M416 5 76 418 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=79310 $D=1
M417 6 76 419 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=83940 $D=1
M418 420 77 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=79310 $D=1
M419 421 77 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=83940 $D=1
M420 422 76 212 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=79310 $D=1
M421 423 76 213 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=83940 $D=1
M422 5 422 730 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=79310 $D=1
M423 6 423 731 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=83940 $D=1
M424 424 730 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=79310 $D=1
M425 425 731 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=83940 $D=1
M426 422 418 424 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=79310 $D=1
M427 423 419 425 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=83940 $D=1
M428 424 77 222 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=79310 $D=1
M429 425 77 223 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=83940 $D=1
M430 226 78 424 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=79310 $D=1
M431 227 78 425 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=83940 $D=1
M432 426 78 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=79310 $D=1
M433 427 78 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=83940 $D=1
M434 5 79 428 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=79310 $D=1
M435 6 79 429 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=83940 $D=1
M436 430 80 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=79310 $D=1
M437 431 80 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=83940 $D=1
M438 432 79 212 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=79310 $D=1
M439 433 79 213 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=83940 $D=1
M440 5 432 732 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=79310 $D=1
M441 6 433 733 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=83940 $D=1
M442 434 732 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=79310 $D=1
M443 435 733 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=83940 $D=1
M444 432 428 434 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=79310 $D=1
M445 433 429 435 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=83940 $D=1
M446 434 80 222 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=79310 $D=1
M447 435 80 223 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=83940 $D=1
M448 226 81 434 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=79310 $D=1
M449 227 81 435 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=83940 $D=1
M450 436 81 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=79310 $D=1
M451 437 81 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=83940 $D=1
M452 5 82 438 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=79310 $D=1
M453 6 82 439 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=83940 $D=1
M454 440 83 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=79310 $D=1
M455 441 83 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=83940 $D=1
M456 442 82 212 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=79310 $D=1
M457 443 82 213 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=83940 $D=1
M458 5 442 734 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=79310 $D=1
M459 6 443 735 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=83940 $D=1
M460 444 734 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=79310 $D=1
M461 445 735 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=83940 $D=1
M462 442 438 444 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=79310 $D=1
M463 443 439 445 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=83940 $D=1
M464 444 83 222 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=79310 $D=1
M465 445 83 223 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=83940 $D=1
M466 226 84 444 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=79310 $D=1
M467 227 84 445 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=83940 $D=1
M468 446 84 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=79310 $D=1
M469 447 84 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=83940 $D=1
M470 5 85 448 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=79310 $D=1
M471 6 85 449 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=83940 $D=1
M472 450 86 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=79310 $D=1
M473 451 86 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=83940 $D=1
M474 452 85 212 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=79310 $D=1
M475 453 85 213 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=83940 $D=1
M476 5 452 736 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=79310 $D=1
M477 6 453 737 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=83940 $D=1
M478 454 736 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=79310 $D=1
M479 455 737 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=83940 $D=1
M480 452 448 454 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=79310 $D=1
M481 453 449 455 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=83940 $D=1
M482 454 86 222 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=79310 $D=1
M483 455 86 223 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=83940 $D=1
M484 226 87 454 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=79310 $D=1
M485 227 87 455 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=83940 $D=1
M486 456 87 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=79310 $D=1
M487 457 87 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=83940 $D=1
M488 5 88 458 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=79310 $D=1
M489 6 88 459 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=83940 $D=1
M490 460 89 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=79310 $D=1
M491 461 89 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=83940 $D=1
M492 462 88 212 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=79310 $D=1
M493 463 88 213 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=83940 $D=1
M494 5 462 738 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=79310 $D=1
M495 6 463 739 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=83940 $D=1
M496 464 738 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=79310 $D=1
M497 465 739 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=83940 $D=1
M498 462 458 464 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=79310 $D=1
M499 463 459 465 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=83940 $D=1
M500 464 89 222 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=79310 $D=1
M501 465 89 223 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=83940 $D=1
M502 226 90 464 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=79310 $D=1
M503 227 90 465 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=83940 $D=1
M504 466 90 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=79310 $D=1
M505 467 90 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=83940 $D=1
M506 5 91 468 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=79310 $D=1
M507 6 91 469 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=83940 $D=1
M508 470 92 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=79310 $D=1
M509 471 92 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=83940 $D=1
M510 472 91 212 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=79310 $D=1
M511 473 91 213 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=83940 $D=1
M512 5 472 740 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=79310 $D=1
M513 6 473 741 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=83940 $D=1
M514 474 740 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=79310 $D=1
M515 475 741 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=83940 $D=1
M516 472 468 474 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=79310 $D=1
M517 473 469 475 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=83940 $D=1
M518 474 92 222 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=79310 $D=1
M519 475 92 223 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=83940 $D=1
M520 226 93 474 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=79310 $D=1
M521 227 93 475 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=83940 $D=1
M522 476 93 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=79310 $D=1
M523 477 93 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=83940 $D=1
M524 5 94 478 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=79310 $D=1
M525 6 94 479 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=83940 $D=1
M526 480 95 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=79310 $D=1
M527 481 95 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=83940 $D=1
M528 482 94 212 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=79310 $D=1
M529 483 94 213 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=83940 $D=1
M530 5 482 742 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=79310 $D=1
M531 6 483 743 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=83940 $D=1
M532 484 742 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=79310 $D=1
M533 485 743 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=83940 $D=1
M534 482 478 484 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=79310 $D=1
M535 483 479 485 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=83940 $D=1
M536 484 95 222 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=79310 $D=1
M537 485 95 223 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=83940 $D=1
M538 226 96 484 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=79310 $D=1
M539 227 96 485 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=83940 $D=1
M540 486 96 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=79310 $D=1
M541 487 96 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=83940 $D=1
M542 5 97 488 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=79310 $D=1
M543 6 97 489 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=83940 $D=1
M544 490 98 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=79310 $D=1
M545 491 98 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=83940 $D=1
M546 492 97 212 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=79310 $D=1
M547 493 97 213 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=83940 $D=1
M548 5 492 744 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=79310 $D=1
M549 6 493 745 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=83940 $D=1
M550 494 744 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=79310 $D=1
M551 495 745 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=83940 $D=1
M552 492 488 494 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=79310 $D=1
M553 493 489 495 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=83940 $D=1
M554 494 98 222 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=79310 $D=1
M555 495 98 223 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=83940 $D=1
M556 226 99 494 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=79310 $D=1
M557 227 99 495 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=83940 $D=1
M558 496 99 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=79310 $D=1
M559 497 99 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=83940 $D=1
M560 5 100 498 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=79310 $D=1
M561 6 100 499 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=83940 $D=1
M562 500 101 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=79310 $D=1
M563 501 101 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=83940 $D=1
M564 502 100 212 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=79310 $D=1
M565 503 100 213 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=83940 $D=1
M566 5 502 746 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=79310 $D=1
M567 6 503 747 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=83940 $D=1
M568 504 746 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=79310 $D=1
M569 505 747 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=83940 $D=1
M570 502 498 504 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=79310 $D=1
M571 503 499 505 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=83940 $D=1
M572 504 101 222 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=79310 $D=1
M573 505 101 223 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=83940 $D=1
M574 226 102 504 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=79310 $D=1
M575 227 102 505 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=83940 $D=1
M576 506 102 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=79310 $D=1
M577 507 102 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=83940 $D=1
M578 5 103 508 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=79310 $D=1
M579 6 103 509 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=83940 $D=1
M580 510 104 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=79310 $D=1
M581 511 104 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=83940 $D=1
M582 512 103 212 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=79310 $D=1
M583 513 103 213 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=83940 $D=1
M584 5 512 748 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=79310 $D=1
M585 6 513 749 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=83940 $D=1
M586 514 748 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=79310 $D=1
M587 515 749 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=83940 $D=1
M588 512 508 514 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=79310 $D=1
M589 513 509 515 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=83940 $D=1
M590 514 104 222 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=79310 $D=1
M591 515 104 223 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=83940 $D=1
M592 226 105 514 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=79310 $D=1
M593 227 105 515 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=83940 $D=1
M594 516 105 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=79310 $D=1
M595 517 105 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=83940 $D=1
M596 5 106 518 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=79310 $D=1
M597 6 106 519 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=83940 $D=1
M598 520 107 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=79310 $D=1
M599 521 107 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=83940 $D=1
M600 522 106 212 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=79310 $D=1
M601 523 106 213 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=83940 $D=1
M602 5 522 750 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=79310 $D=1
M603 6 523 751 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=83940 $D=1
M604 524 750 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=79310 $D=1
M605 525 751 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=83940 $D=1
M606 522 518 524 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=79310 $D=1
M607 523 519 525 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=83940 $D=1
M608 524 107 222 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=79310 $D=1
M609 525 107 223 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=83940 $D=1
M610 226 108 524 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=79310 $D=1
M611 227 108 525 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=83940 $D=1
M612 526 108 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=79310 $D=1
M613 527 108 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=83940 $D=1
M614 5 109 528 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=79310 $D=1
M615 6 109 529 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=83940 $D=1
M616 530 110 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=79310 $D=1
M617 531 110 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=83940 $D=1
M618 5 110 222 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=79310 $D=1
M619 6 110 223 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=83940 $D=1
M620 226 109 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=79310 $D=1
M621 227 109 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=83940 $D=1
M622 5 534 532 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=79310 $D=1
M623 6 535 533 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=83940 $D=1
M624 534 111 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=79310 $D=1
M625 535 111 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=83940 $D=1
M626 752 222 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=79310 $D=1
M627 753 223 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=83940 $D=1
M628 536 532 752 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=79310 $D=1
M629 537 533 753 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=83940 $D=1
M630 5 536 538 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=79310 $D=1
M631 6 537 539 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=83940 $D=1
M632 754 538 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=79310 $D=1
M633 755 539 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=83940 $D=1
M634 536 534 754 5 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=79310 $D=1
M635 537 535 755 6 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=83940 $D=1
M636 5 542 540 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=79310 $D=1
M637 6 543 541 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=83940 $D=1
M638 542 111 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=79310 $D=1
M639 543 111 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=83940 $D=1
M640 756 226 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=79310 $D=1
M641 757 227 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=83940 $D=1
M642 544 540 756 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=79310 $D=1
M643 545 541 757 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=83940 $D=1
M644 5 544 112 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=79310 $D=1
M645 6 545 113 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=83940 $D=1
M646 758 112 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=79310 $D=1
M647 759 113 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=83940 $D=1
M648 544 542 758 5 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=79310 $D=1
M649 545 543 759 6 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=83940 $D=1
M650 546 114 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=79310 $D=1
M651 547 114 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=83940 $D=1
M652 548 546 538 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=79310 $D=1
M653 549 547 539 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=83940 $D=1
M654 115 114 548 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=79310 $D=1
M655 116 114 549 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=83940 $D=1
M656 550 117 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=79310 $D=1
M657 551 117 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=83940 $D=1
M658 552 550 112 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=79310 $D=1
M659 553 551 113 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=83940 $D=1
M660 760 117 552 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=79310 $D=1
M661 761 117 553 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=83940 $D=1
M662 5 112 760 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=79310 $D=1
M663 6 113 761 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=83940 $D=1
M664 554 118 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=79310 $D=1
M665 555 118 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=83940 $D=1
M666 556 554 552 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=79310 $D=1
M667 557 555 553 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=83940 $D=1
M668 10 118 556 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=79310 $D=1
M669 11 118 557 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=83940 $D=1
M670 559 558 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=79310 $D=1
M671 560 119 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=83940 $D=1
M672 5 563 561 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=79310 $D=1
M673 6 564 562 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=83940 $D=1
M674 565 548 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=79310 $D=1
M675 566 549 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=83940 $D=1
M676 563 565 558 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=79310 $D=1
M677 564 566 119 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=83940 $D=1
M678 559 548 563 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=79310 $D=1
M679 560 549 564 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=83940 $D=1
M680 567 561 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=79310 $D=1
M681 568 562 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=83940 $D=1
M682 120 567 556 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=79310 $D=1
M683 558 568 557 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=83940 $D=1
M684 548 561 120 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=79310 $D=1
M685 549 562 558 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=83940 $D=1
M686 569 120 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=79310 $D=1
M687 570 558 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=83940 $D=1
M688 571 561 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=79310 $D=1
M689 572 562 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=83940 $D=1
M690 573 571 569 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=79310 $D=1
M691 574 572 570 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=83940 $D=1
M692 556 561 573 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=79310 $D=1
M693 557 562 574 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=83940 $D=1
M694 575 548 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=79310 $D=1
M695 576 549 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=83940 $D=1
M696 5 556 575 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=79310 $D=1
M697 6 557 576 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=83940 $D=1
M698 577 573 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=79310 $D=1
M699 578 574 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=83940 $D=1
M700 790 548 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=79310 $D=1
M701 791 549 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=83940 $D=1
M702 579 556 790 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=79310 $D=1
M703 580 557 791 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=83940 $D=1
M704 792 548 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=79310 $D=1
M705 793 549 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=83940 $D=1
M706 581 556 792 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=79310 $D=1
M707 582 557 793 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=83940 $D=1
M708 585 548 583 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=79310 $D=1
M709 586 549 584 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=83940 $D=1
M710 583 556 585 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=79310 $D=1
M711 584 557 586 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=83940 $D=1
M712 5 581 583 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=79310 $D=1
M713 6 582 584 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=83940 $D=1
M714 587 123 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=79310 $D=1
M715 588 123 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=83940 $D=1
M716 589 587 575 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=79310 $D=1
M717 590 588 576 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=83940 $D=1
M718 579 123 589 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=79310 $D=1
M719 580 123 590 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=83940 $D=1
M720 591 587 577 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=79310 $D=1
M721 592 588 578 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=83940 $D=1
M722 585 123 591 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=79310 $D=1
M723 586 123 592 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=83940 $D=1
M724 593 124 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=79310 $D=1
M725 594 124 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=83940 $D=1
M726 595 593 591 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=79310 $D=1
M727 596 594 592 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=83940 $D=1
M728 589 124 595 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=79310 $D=1
M729 590 124 596 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=83940 $D=1
M730 12 595 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=79310 $D=1
M731 13 596 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=83940 $D=1
M732 597 125 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=79310 $D=1
M733 598 125 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=83940 $D=1
M734 599 597 126 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=79310 $D=1
M735 600 598 127 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=83940 $D=1
M736 128 125 599 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=79310 $D=1
M737 129 125 600 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=83940 $D=1
M738 601 125 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=79310 $D=1
M739 602 125 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=83940 $D=1
M740 606 601 130 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=79310 $D=1
M741 607 602 132 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=83940 $D=1
M742 133 125 606 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=79310 $D=1
M743 131 125 607 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=83940 $D=1
M744 608 125 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=79310 $D=1
M745 609 125 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=83940 $D=1
M746 610 608 134 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=79310 $D=1
M747 611 609 135 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=83940 $D=1
M748 136 125 610 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=79310 $D=1
M749 137 125 611 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=83940 $D=1
M750 612 125 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=79310 $D=1
M751 613 125 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=83940 $D=1
M752 614 612 138 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=79310 $D=1
M753 615 613 139 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=83940 $D=1
M754 140 125 614 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=79310 $D=1
M755 141 125 615 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=83940 $D=1
M756 616 125 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=79310 $D=1
M757 617 125 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=83940 $D=1
M758 618 616 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=79310 $D=1
M759 619 617 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=83940 $D=1
M760 142 125 618 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=79310 $D=1
M761 143 125 619 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=83940 $D=1
M762 5 548 772 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=79310 $D=1
M763 6 549 773 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=83940 $D=1
M764 129 772 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=79310 $D=1
M765 126 773 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=83940 $D=1
M766 620 144 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=79310 $D=1
M767 621 144 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=83940 $D=1
M768 145 620 129 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=79310 $D=1
M769 146 621 126 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=83940 $D=1
M770 599 144 145 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=79310 $D=1
M771 600 144 146 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=83940 $D=1
M772 622 147 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=79310 $D=1
M773 623 147 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=83940 $D=1
M774 122 622 145 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=79310 $D=1
M775 121 623 146 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=83940 $D=1
M776 606 147 122 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=79310 $D=1
M777 607 147 121 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=83940 $D=1
M778 624 148 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=79310 $D=1
M779 625 148 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=83940 $D=1
M780 149 624 122 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=79310 $D=1
M781 150 625 121 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=83940 $D=1
M782 610 148 149 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=79310 $D=1
M783 611 148 150 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=83940 $D=1
M784 626 151 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=79310 $D=1
M785 627 151 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=83940 $D=1
M786 152 626 149 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=79310 $D=1
M787 153 627 150 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=83940 $D=1
M788 614 151 152 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=79310 $D=1
M789 615 151 153 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=83940 $D=1
M790 628 154 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=79310 $D=1
M791 629 154 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=83940 $D=1
M792 198 628 152 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=79310 $D=1
M793 199 629 153 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=83940 $D=1
M794 618 154 198 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=79310 $D=1
M795 619 154 199 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=83940 $D=1
M796 630 155 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=79310 $D=1
M797 631 155 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=83940 $D=1
M798 632 630 112 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=79310 $D=1
M799 633 631 113 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=83940 $D=1
M800 10 155 632 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=79310 $D=1
M801 11 155 633 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=83940 $D=1
M802 794 538 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=79310 $D=1
M803 795 539 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=83940 $D=1
M804 634 632 794 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=79310 $D=1
M805 635 633 795 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=83940 $D=1
M806 638 538 636 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=79310 $D=1
M807 639 539 637 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=83940 $D=1
M808 636 632 638 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=79310 $D=1
M809 637 633 639 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=83940 $D=1
M810 5 634 636 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=79310 $D=1
M811 6 635 637 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=83940 $D=1
M812 796 640 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=79310 $D=1
M813 797 641 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=83940 $D=1
M814 774 638 796 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=79310 $D=1
M815 775 639 797 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=83940 $D=1
M816 641 774 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=79310 $D=1
M817 156 775 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=83940 $D=1
M818 642 538 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=79310 $D=1
M819 643 539 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=83940 $D=1
M820 5 644 642 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=79310 $D=1
M821 6 645 643 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=83940 $D=1
M822 644 632 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=79310 $D=1
M823 645 633 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=83940 $D=1
M824 798 642 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=79310 $D=1
M825 799 643 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=83940 $D=1
M826 646 640 798 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=79310 $D=1
M827 647 641 799 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=83940 $D=1
M828 649 157 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=79310 $D=1
M829 650 648 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=83940 $D=1
M830 800 646 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=79310 $D=1
M831 801 647 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=83940 $D=1
M832 648 649 800 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=79310 $D=1
M833 158 650 801 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=83940 $D=1
M834 652 651 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=79310 $D=1
M835 653 159 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=83940 $D=1
M836 5 656 654 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=79310 $D=1
M837 6 657 655 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=83940 $D=1
M838 658 115 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=79310 $D=1
M839 659 116 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=83940 $D=1
M840 656 658 651 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=79310 $D=1
M841 657 659 159 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=83940 $D=1
M842 652 115 656 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=79310 $D=1
M843 653 116 657 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=83940 $D=1
M844 660 654 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=79310 $D=1
M845 661 655 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=83940 $D=1
M846 160 660 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=79310 $D=1
M847 651 661 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=83940 $D=1
M848 115 654 160 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=79310 $D=1
M849 116 655 651 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=83940 $D=1
M850 662 160 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=79310 $D=1
M851 663 651 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=83940 $D=1
M852 664 654 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=79310 $D=1
M853 665 655 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=83940 $D=1
M854 200 664 662 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=79310 $D=1
M855 201 665 663 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=83940 $D=1
M856 5 654 200 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=79310 $D=1
M857 6 655 201 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=83940 $D=1
M858 666 161 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=79310 $D=1
M859 667 161 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=83940 $D=1
M860 668 666 200 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=79310 $D=1
M861 669 667 201 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=83940 $D=1
M862 12 161 668 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=79310 $D=1
M863 13 161 669 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=83940 $D=1
M864 670 162 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=79310 $D=1
M865 671 162 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=83940 $D=1
M866 162 670 668 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=79310 $D=1
M867 162 671 669 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=83940 $D=1
M868 5 162 162 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=79310 $D=1
M869 6 162 162 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=83940 $D=1
M870 672 111 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=79310 $D=1
M871 673 111 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=83940 $D=1
M872 5 672 674 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=79310 $D=1
M873 6 673 675 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=83940 $D=1
M874 676 111 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=79310 $D=1
M875 677 111 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=83940 $D=1
M876 678 672 162 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=79310 $D=1
M877 679 673 162 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=83940 $D=1
M878 5 678 776 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=79310 $D=1
M879 6 679 777 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=83940 $D=1
M880 680 776 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=79310 $D=1
M881 681 777 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=83940 $D=1
M882 678 674 680 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=79310 $D=1
M883 679 675 681 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=83940 $D=1
M884 682 111 680 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=79310 $D=1
M885 683 111 681 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=83940 $D=1
M886 5 686 684 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=79310 $D=1
M887 6 687 685 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=83940 $D=1
M888 686 111 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=79310 $D=1
M889 687 111 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=83940 $D=1
M890 778 682 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=79310 $D=1
M891 779 683 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=83940 $D=1
M892 688 684 778 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=79310 $D=1
M893 689 685 779 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=83940 $D=1
M894 5 688 115 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=79310 $D=1
M895 6 689 116 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=83940 $D=1
M896 780 115 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=79310 $D=1
M897 781 116 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=83940 $D=1
M898 688 686 780 5 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=79310 $D=1
M899 689 687 781 6 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=83940 $D=1
M900 174 1 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=80560 $D=0
M901 175 1 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=85190 $D=0
M902 176 1 2 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=80560 $D=0
M903 177 1 3 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=85190 $D=0
M904 5 174 176 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=80560 $D=0
M905 6 175 177 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=85190 $D=0
M906 178 1 4 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=80560 $D=0
M907 179 1 4 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=85190 $D=0
M908 2 174 178 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=80560 $D=0
M909 3 175 179 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=85190 $D=0
M910 180 1 5 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=80560 $D=0
M911 181 1 6 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=85190 $D=0
M912 2 174 180 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=80560 $D=0
M913 3 175 181 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=85190 $D=0
M914 184 7 180 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=80560 $D=0
M915 185 7 181 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=85190 $D=0
M916 182 7 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=80560 $D=0
M917 183 7 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=85190 $D=0
M918 186 7 178 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=80560 $D=0
M919 187 7 179 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=85190 $D=0
M920 176 182 186 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=80560 $D=0
M921 177 183 187 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=85190 $D=0
M922 188 8 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=80560 $D=0
M923 189 8 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=85190 $D=0
M924 190 8 186 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=80560 $D=0
M925 191 8 187 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=85190 $D=0
M926 184 188 190 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=80560 $D=0
M927 185 189 191 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=85190 $D=0
M928 192 9 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=80560 $D=0
M929 193 9 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=85190 $D=0
M930 194 9 5 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=80560 $D=0
M931 195 9 6 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=85190 $D=0
M932 10 192 194 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=80560 $D=0
M933 11 193 195 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=85190 $D=0
M934 196 9 12 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=80560 $D=0
M935 197 9 13 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=85190 $D=0
M936 198 192 196 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=80560 $D=0
M937 199 193 197 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=85190 $D=0
M938 202 9 200 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=80560 $D=0
M939 203 9 201 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=85190 $D=0
M940 190 192 202 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=80560 $D=0
M941 191 193 203 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=85190 $D=0
M942 206 14 202 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=80560 $D=0
M943 207 14 203 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=85190 $D=0
M944 204 14 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=80560 $D=0
M945 205 14 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=85190 $D=0
M946 208 14 196 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=80560 $D=0
M947 209 14 197 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=85190 $D=0
M948 194 204 208 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=80560 $D=0
M949 195 205 209 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=85190 $D=0
M950 210 15 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=80560 $D=0
M951 211 15 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=85190 $D=0
M952 212 15 208 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=80560 $D=0
M953 213 15 209 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=85190 $D=0
M954 206 210 212 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=80560 $D=0
M955 207 211 213 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=85190 $D=0
M956 163 16 214 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=80560 $D=0
M957 164 16 215 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=85190 $D=0
M958 216 17 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=80560 $D=0
M959 217 17 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=85190 $D=0
M960 218 214 212 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=80560 $D=0
M961 219 215 213 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=85190 $D=0
M962 163 218 690 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=80560 $D=0
M963 164 219 691 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=85190 $D=0
M964 220 690 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=80560 $D=0
M965 221 691 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=85190 $D=0
M966 218 16 220 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=80560 $D=0
M967 219 16 221 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=85190 $D=0
M968 220 216 222 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=80560 $D=0
M969 221 217 223 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=85190 $D=0
M970 226 224 220 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=80560 $D=0
M971 227 225 221 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=85190 $D=0
M972 224 18 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=80560 $D=0
M973 225 18 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=85190 $D=0
M974 163 19 228 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=80560 $D=0
M975 164 19 229 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=85190 $D=0
M976 230 20 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=80560 $D=0
M977 231 20 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=85190 $D=0
M978 232 228 212 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=80560 $D=0
M979 233 229 213 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=85190 $D=0
M980 163 232 692 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=80560 $D=0
M981 164 233 693 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=85190 $D=0
M982 234 692 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=80560 $D=0
M983 235 693 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=85190 $D=0
M984 232 19 234 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=80560 $D=0
M985 233 19 235 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=85190 $D=0
M986 234 230 222 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=80560 $D=0
M987 235 231 223 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=85190 $D=0
M988 226 236 234 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=80560 $D=0
M989 227 237 235 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=85190 $D=0
M990 236 21 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=80560 $D=0
M991 237 21 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=85190 $D=0
M992 163 22 238 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=80560 $D=0
M993 164 22 239 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=85190 $D=0
M994 240 23 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=80560 $D=0
M995 241 23 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=85190 $D=0
M996 242 238 212 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=80560 $D=0
M997 243 239 213 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=85190 $D=0
M998 163 242 694 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=80560 $D=0
M999 164 243 695 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=85190 $D=0
M1000 244 694 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=80560 $D=0
M1001 245 695 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=85190 $D=0
M1002 242 22 244 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=80560 $D=0
M1003 243 22 245 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=85190 $D=0
M1004 244 240 222 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=80560 $D=0
M1005 245 241 223 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=85190 $D=0
M1006 226 246 244 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=80560 $D=0
M1007 227 247 245 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=85190 $D=0
M1008 246 24 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=80560 $D=0
M1009 247 24 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=85190 $D=0
M1010 163 25 248 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=80560 $D=0
M1011 164 25 249 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=85190 $D=0
M1012 250 26 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=80560 $D=0
M1013 251 26 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=85190 $D=0
M1014 252 248 212 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=80560 $D=0
M1015 253 249 213 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=85190 $D=0
M1016 163 252 696 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=80560 $D=0
M1017 164 253 697 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=85190 $D=0
M1018 254 696 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=80560 $D=0
M1019 255 697 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=85190 $D=0
M1020 252 25 254 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=80560 $D=0
M1021 253 25 255 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=85190 $D=0
M1022 254 250 222 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=80560 $D=0
M1023 255 251 223 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=85190 $D=0
M1024 226 256 254 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=80560 $D=0
M1025 227 257 255 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=85190 $D=0
M1026 256 27 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=80560 $D=0
M1027 257 27 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=85190 $D=0
M1028 163 28 258 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=80560 $D=0
M1029 164 28 259 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=85190 $D=0
M1030 260 29 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=80560 $D=0
M1031 261 29 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=85190 $D=0
M1032 262 258 212 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=80560 $D=0
M1033 263 259 213 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=85190 $D=0
M1034 163 262 698 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=80560 $D=0
M1035 164 263 699 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=85190 $D=0
M1036 264 698 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=80560 $D=0
M1037 265 699 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=85190 $D=0
M1038 262 28 264 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=80560 $D=0
M1039 263 28 265 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=85190 $D=0
M1040 264 260 222 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=80560 $D=0
M1041 265 261 223 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=85190 $D=0
M1042 226 266 264 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=80560 $D=0
M1043 227 267 265 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=85190 $D=0
M1044 266 30 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=80560 $D=0
M1045 267 30 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=85190 $D=0
M1046 163 31 268 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=80560 $D=0
M1047 164 31 269 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=85190 $D=0
M1048 270 32 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=80560 $D=0
M1049 271 32 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=85190 $D=0
M1050 272 268 212 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=80560 $D=0
M1051 273 269 213 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=85190 $D=0
M1052 163 272 700 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=80560 $D=0
M1053 164 273 701 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=85190 $D=0
M1054 274 700 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=80560 $D=0
M1055 275 701 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=85190 $D=0
M1056 272 31 274 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=80560 $D=0
M1057 273 31 275 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=85190 $D=0
M1058 274 270 222 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=80560 $D=0
M1059 275 271 223 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=85190 $D=0
M1060 226 276 274 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=80560 $D=0
M1061 227 277 275 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=85190 $D=0
M1062 276 33 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=80560 $D=0
M1063 277 33 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=85190 $D=0
M1064 163 34 278 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=80560 $D=0
M1065 164 34 279 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=85190 $D=0
M1066 280 35 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=80560 $D=0
M1067 281 35 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=85190 $D=0
M1068 282 278 212 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=80560 $D=0
M1069 283 279 213 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=85190 $D=0
M1070 163 282 702 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=80560 $D=0
M1071 164 283 703 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=85190 $D=0
M1072 284 702 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=80560 $D=0
M1073 285 703 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=85190 $D=0
M1074 282 34 284 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=80560 $D=0
M1075 283 34 285 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=85190 $D=0
M1076 284 280 222 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=80560 $D=0
M1077 285 281 223 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=85190 $D=0
M1078 226 286 284 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=80560 $D=0
M1079 227 287 285 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=85190 $D=0
M1080 286 36 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=80560 $D=0
M1081 287 36 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=85190 $D=0
M1082 163 37 288 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=80560 $D=0
M1083 164 37 289 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=85190 $D=0
M1084 290 38 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=80560 $D=0
M1085 291 38 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=85190 $D=0
M1086 292 288 212 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=80560 $D=0
M1087 293 289 213 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=85190 $D=0
M1088 163 292 704 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=80560 $D=0
M1089 164 293 705 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=85190 $D=0
M1090 294 704 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=80560 $D=0
M1091 295 705 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=85190 $D=0
M1092 292 37 294 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=80560 $D=0
M1093 293 37 295 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=85190 $D=0
M1094 294 290 222 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=80560 $D=0
M1095 295 291 223 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=85190 $D=0
M1096 226 296 294 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=80560 $D=0
M1097 227 297 295 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=85190 $D=0
M1098 296 39 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=80560 $D=0
M1099 297 39 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=85190 $D=0
M1100 163 40 298 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=80560 $D=0
M1101 164 40 299 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=85190 $D=0
M1102 300 41 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=80560 $D=0
M1103 301 41 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=85190 $D=0
M1104 302 298 212 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=80560 $D=0
M1105 303 299 213 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=85190 $D=0
M1106 163 302 706 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=80560 $D=0
M1107 164 303 707 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=85190 $D=0
M1108 304 706 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=80560 $D=0
M1109 305 707 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=85190 $D=0
M1110 302 40 304 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=80560 $D=0
M1111 303 40 305 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=85190 $D=0
M1112 304 300 222 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=80560 $D=0
M1113 305 301 223 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=85190 $D=0
M1114 226 306 304 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=80560 $D=0
M1115 227 307 305 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=85190 $D=0
M1116 306 42 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=80560 $D=0
M1117 307 42 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=85190 $D=0
M1118 163 43 308 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=80560 $D=0
M1119 164 43 309 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=85190 $D=0
M1120 310 44 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=80560 $D=0
M1121 311 44 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=85190 $D=0
M1122 312 308 212 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=80560 $D=0
M1123 313 309 213 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=85190 $D=0
M1124 163 312 708 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=80560 $D=0
M1125 164 313 709 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=85190 $D=0
M1126 314 708 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=80560 $D=0
M1127 315 709 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=85190 $D=0
M1128 312 43 314 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=80560 $D=0
M1129 313 43 315 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=85190 $D=0
M1130 314 310 222 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=80560 $D=0
M1131 315 311 223 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=85190 $D=0
M1132 226 316 314 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=80560 $D=0
M1133 227 317 315 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=85190 $D=0
M1134 316 45 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=80560 $D=0
M1135 317 45 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=85190 $D=0
M1136 163 46 318 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=80560 $D=0
M1137 164 46 319 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=85190 $D=0
M1138 320 47 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=80560 $D=0
M1139 321 47 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=85190 $D=0
M1140 322 318 212 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=80560 $D=0
M1141 323 319 213 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=85190 $D=0
M1142 163 322 710 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=80560 $D=0
M1143 164 323 711 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=85190 $D=0
M1144 324 710 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=80560 $D=0
M1145 325 711 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=85190 $D=0
M1146 322 46 324 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=80560 $D=0
M1147 323 46 325 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=85190 $D=0
M1148 324 320 222 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=80560 $D=0
M1149 325 321 223 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=85190 $D=0
M1150 226 326 324 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=80560 $D=0
M1151 227 327 325 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=85190 $D=0
M1152 326 48 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=80560 $D=0
M1153 327 48 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=85190 $D=0
M1154 163 49 328 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=80560 $D=0
M1155 164 49 329 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=85190 $D=0
M1156 330 50 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=80560 $D=0
M1157 331 50 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=85190 $D=0
M1158 332 328 212 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=80560 $D=0
M1159 333 329 213 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=85190 $D=0
M1160 163 332 712 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=80560 $D=0
M1161 164 333 713 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=85190 $D=0
M1162 334 712 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=80560 $D=0
M1163 335 713 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=85190 $D=0
M1164 332 49 334 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=80560 $D=0
M1165 333 49 335 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=85190 $D=0
M1166 334 330 222 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=80560 $D=0
M1167 335 331 223 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=85190 $D=0
M1168 226 336 334 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=80560 $D=0
M1169 227 337 335 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=85190 $D=0
M1170 336 51 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=80560 $D=0
M1171 337 51 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=85190 $D=0
M1172 163 52 338 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=80560 $D=0
M1173 164 52 339 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=85190 $D=0
M1174 340 53 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=80560 $D=0
M1175 341 53 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=85190 $D=0
M1176 342 338 212 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=80560 $D=0
M1177 343 339 213 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=85190 $D=0
M1178 163 342 714 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=80560 $D=0
M1179 164 343 715 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=85190 $D=0
M1180 344 714 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=80560 $D=0
M1181 345 715 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=85190 $D=0
M1182 342 52 344 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=80560 $D=0
M1183 343 52 345 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=85190 $D=0
M1184 344 340 222 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=80560 $D=0
M1185 345 341 223 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=85190 $D=0
M1186 226 346 344 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=80560 $D=0
M1187 227 347 345 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=85190 $D=0
M1188 346 54 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=80560 $D=0
M1189 347 54 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=85190 $D=0
M1190 163 55 348 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=80560 $D=0
M1191 164 55 349 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=85190 $D=0
M1192 350 56 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=80560 $D=0
M1193 351 56 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=85190 $D=0
M1194 352 348 212 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=80560 $D=0
M1195 353 349 213 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=85190 $D=0
M1196 163 352 716 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=80560 $D=0
M1197 164 353 717 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=85190 $D=0
M1198 354 716 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=80560 $D=0
M1199 355 717 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=85190 $D=0
M1200 352 55 354 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=80560 $D=0
M1201 353 55 355 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=85190 $D=0
M1202 354 350 222 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=80560 $D=0
M1203 355 351 223 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=85190 $D=0
M1204 226 356 354 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=80560 $D=0
M1205 227 357 355 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=85190 $D=0
M1206 356 57 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=80560 $D=0
M1207 357 57 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=85190 $D=0
M1208 163 58 358 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=80560 $D=0
M1209 164 58 359 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=85190 $D=0
M1210 360 59 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=80560 $D=0
M1211 361 59 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=85190 $D=0
M1212 362 358 212 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=80560 $D=0
M1213 363 359 213 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=85190 $D=0
M1214 163 362 718 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=80560 $D=0
M1215 164 363 719 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=85190 $D=0
M1216 364 718 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=80560 $D=0
M1217 365 719 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=85190 $D=0
M1218 362 58 364 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=80560 $D=0
M1219 363 58 365 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=85190 $D=0
M1220 364 360 222 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=80560 $D=0
M1221 365 361 223 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=85190 $D=0
M1222 226 366 364 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=80560 $D=0
M1223 227 367 365 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=85190 $D=0
M1224 366 60 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=80560 $D=0
M1225 367 60 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=85190 $D=0
M1226 163 61 368 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=80560 $D=0
M1227 164 61 369 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=85190 $D=0
M1228 370 62 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=80560 $D=0
M1229 371 62 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=85190 $D=0
M1230 372 368 212 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=80560 $D=0
M1231 373 369 213 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=85190 $D=0
M1232 163 372 720 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=80560 $D=0
M1233 164 373 721 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=85190 $D=0
M1234 374 720 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=80560 $D=0
M1235 375 721 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=85190 $D=0
M1236 372 61 374 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=80560 $D=0
M1237 373 61 375 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=85190 $D=0
M1238 374 370 222 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=80560 $D=0
M1239 375 371 223 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=85190 $D=0
M1240 226 376 374 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=80560 $D=0
M1241 227 377 375 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=85190 $D=0
M1242 376 63 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=80560 $D=0
M1243 377 63 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=85190 $D=0
M1244 163 64 378 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=80560 $D=0
M1245 164 64 379 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=85190 $D=0
M1246 380 65 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=80560 $D=0
M1247 381 65 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=85190 $D=0
M1248 382 378 212 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=80560 $D=0
M1249 383 379 213 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=85190 $D=0
M1250 163 382 722 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=80560 $D=0
M1251 164 383 723 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=85190 $D=0
M1252 384 722 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=80560 $D=0
M1253 385 723 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=85190 $D=0
M1254 382 64 384 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=80560 $D=0
M1255 383 64 385 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=85190 $D=0
M1256 384 380 222 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=80560 $D=0
M1257 385 381 223 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=85190 $D=0
M1258 226 386 384 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=80560 $D=0
M1259 227 387 385 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=85190 $D=0
M1260 386 66 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=80560 $D=0
M1261 387 66 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=85190 $D=0
M1262 163 67 388 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=80560 $D=0
M1263 164 67 389 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=85190 $D=0
M1264 390 68 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=80560 $D=0
M1265 391 68 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=85190 $D=0
M1266 392 388 212 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=80560 $D=0
M1267 393 389 213 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=85190 $D=0
M1268 163 392 724 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=80560 $D=0
M1269 164 393 725 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=85190 $D=0
M1270 394 724 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=80560 $D=0
M1271 395 725 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=85190 $D=0
M1272 392 67 394 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=80560 $D=0
M1273 393 67 395 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=85190 $D=0
M1274 394 390 222 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=80560 $D=0
M1275 395 391 223 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=85190 $D=0
M1276 226 396 394 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=80560 $D=0
M1277 227 397 395 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=85190 $D=0
M1278 396 69 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=80560 $D=0
M1279 397 69 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=85190 $D=0
M1280 163 70 398 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=80560 $D=0
M1281 164 70 399 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=85190 $D=0
M1282 400 71 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=80560 $D=0
M1283 401 71 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=85190 $D=0
M1284 402 398 212 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=80560 $D=0
M1285 403 399 213 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=85190 $D=0
M1286 163 402 726 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=80560 $D=0
M1287 164 403 727 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=85190 $D=0
M1288 404 726 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=80560 $D=0
M1289 405 727 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=85190 $D=0
M1290 402 70 404 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=80560 $D=0
M1291 403 70 405 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=85190 $D=0
M1292 404 400 222 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=80560 $D=0
M1293 405 401 223 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=85190 $D=0
M1294 226 406 404 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=80560 $D=0
M1295 227 407 405 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=85190 $D=0
M1296 406 72 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=80560 $D=0
M1297 407 72 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=85190 $D=0
M1298 163 73 408 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=80560 $D=0
M1299 164 73 409 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=85190 $D=0
M1300 410 74 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=80560 $D=0
M1301 411 74 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=85190 $D=0
M1302 412 408 212 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=80560 $D=0
M1303 413 409 213 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=85190 $D=0
M1304 163 412 728 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=80560 $D=0
M1305 164 413 729 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=85190 $D=0
M1306 414 728 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=80560 $D=0
M1307 415 729 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=85190 $D=0
M1308 412 73 414 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=80560 $D=0
M1309 413 73 415 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=85190 $D=0
M1310 414 410 222 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=80560 $D=0
M1311 415 411 223 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=85190 $D=0
M1312 226 416 414 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=80560 $D=0
M1313 227 417 415 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=85190 $D=0
M1314 416 75 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=80560 $D=0
M1315 417 75 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=85190 $D=0
M1316 163 76 418 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=80560 $D=0
M1317 164 76 419 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=85190 $D=0
M1318 420 77 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=80560 $D=0
M1319 421 77 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=85190 $D=0
M1320 422 418 212 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=80560 $D=0
M1321 423 419 213 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=85190 $D=0
M1322 163 422 730 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=80560 $D=0
M1323 164 423 731 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=85190 $D=0
M1324 424 730 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=80560 $D=0
M1325 425 731 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=85190 $D=0
M1326 422 76 424 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=80560 $D=0
M1327 423 76 425 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=85190 $D=0
M1328 424 420 222 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=80560 $D=0
M1329 425 421 223 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=85190 $D=0
M1330 226 426 424 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=80560 $D=0
M1331 227 427 425 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=85190 $D=0
M1332 426 78 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=80560 $D=0
M1333 427 78 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=85190 $D=0
M1334 163 79 428 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=80560 $D=0
M1335 164 79 429 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=85190 $D=0
M1336 430 80 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=80560 $D=0
M1337 431 80 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=85190 $D=0
M1338 432 428 212 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=80560 $D=0
M1339 433 429 213 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=85190 $D=0
M1340 163 432 732 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=80560 $D=0
M1341 164 433 733 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=85190 $D=0
M1342 434 732 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=80560 $D=0
M1343 435 733 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=85190 $D=0
M1344 432 79 434 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=80560 $D=0
M1345 433 79 435 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=85190 $D=0
M1346 434 430 222 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=80560 $D=0
M1347 435 431 223 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=85190 $D=0
M1348 226 436 434 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=80560 $D=0
M1349 227 437 435 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=85190 $D=0
M1350 436 81 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=80560 $D=0
M1351 437 81 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=85190 $D=0
M1352 163 82 438 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=80560 $D=0
M1353 164 82 439 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=85190 $D=0
M1354 440 83 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=80560 $D=0
M1355 441 83 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=85190 $D=0
M1356 442 438 212 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=80560 $D=0
M1357 443 439 213 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=85190 $D=0
M1358 163 442 734 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=80560 $D=0
M1359 164 443 735 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=85190 $D=0
M1360 444 734 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=80560 $D=0
M1361 445 735 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=85190 $D=0
M1362 442 82 444 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=80560 $D=0
M1363 443 82 445 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=85190 $D=0
M1364 444 440 222 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=80560 $D=0
M1365 445 441 223 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=85190 $D=0
M1366 226 446 444 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=80560 $D=0
M1367 227 447 445 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=85190 $D=0
M1368 446 84 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=80560 $D=0
M1369 447 84 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=85190 $D=0
M1370 163 85 448 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=80560 $D=0
M1371 164 85 449 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=85190 $D=0
M1372 450 86 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=80560 $D=0
M1373 451 86 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=85190 $D=0
M1374 452 448 212 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=80560 $D=0
M1375 453 449 213 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=85190 $D=0
M1376 163 452 736 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=80560 $D=0
M1377 164 453 737 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=85190 $D=0
M1378 454 736 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=80560 $D=0
M1379 455 737 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=85190 $D=0
M1380 452 85 454 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=80560 $D=0
M1381 453 85 455 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=85190 $D=0
M1382 454 450 222 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=80560 $D=0
M1383 455 451 223 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=85190 $D=0
M1384 226 456 454 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=80560 $D=0
M1385 227 457 455 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=85190 $D=0
M1386 456 87 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=80560 $D=0
M1387 457 87 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=85190 $D=0
M1388 163 88 458 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=80560 $D=0
M1389 164 88 459 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=85190 $D=0
M1390 460 89 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=80560 $D=0
M1391 461 89 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=85190 $D=0
M1392 462 458 212 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=80560 $D=0
M1393 463 459 213 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=85190 $D=0
M1394 163 462 738 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=80560 $D=0
M1395 164 463 739 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=85190 $D=0
M1396 464 738 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=80560 $D=0
M1397 465 739 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=85190 $D=0
M1398 462 88 464 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=80560 $D=0
M1399 463 88 465 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=85190 $D=0
M1400 464 460 222 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=80560 $D=0
M1401 465 461 223 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=85190 $D=0
M1402 226 466 464 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=80560 $D=0
M1403 227 467 465 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=85190 $D=0
M1404 466 90 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=80560 $D=0
M1405 467 90 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=85190 $D=0
M1406 163 91 468 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=80560 $D=0
M1407 164 91 469 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=85190 $D=0
M1408 470 92 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=80560 $D=0
M1409 471 92 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=85190 $D=0
M1410 472 468 212 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=80560 $D=0
M1411 473 469 213 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=85190 $D=0
M1412 163 472 740 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=80560 $D=0
M1413 164 473 741 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=85190 $D=0
M1414 474 740 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=80560 $D=0
M1415 475 741 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=85190 $D=0
M1416 472 91 474 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=80560 $D=0
M1417 473 91 475 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=85190 $D=0
M1418 474 470 222 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=80560 $D=0
M1419 475 471 223 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=85190 $D=0
M1420 226 476 474 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=80560 $D=0
M1421 227 477 475 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=85190 $D=0
M1422 476 93 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=80560 $D=0
M1423 477 93 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=85190 $D=0
M1424 163 94 478 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=80560 $D=0
M1425 164 94 479 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=85190 $D=0
M1426 480 95 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=80560 $D=0
M1427 481 95 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=85190 $D=0
M1428 482 478 212 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=80560 $D=0
M1429 483 479 213 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=85190 $D=0
M1430 163 482 742 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=80560 $D=0
M1431 164 483 743 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=85190 $D=0
M1432 484 742 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=80560 $D=0
M1433 485 743 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=85190 $D=0
M1434 482 94 484 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=80560 $D=0
M1435 483 94 485 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=85190 $D=0
M1436 484 480 222 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=80560 $D=0
M1437 485 481 223 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=85190 $D=0
M1438 226 486 484 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=80560 $D=0
M1439 227 487 485 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=85190 $D=0
M1440 486 96 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=80560 $D=0
M1441 487 96 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=85190 $D=0
M1442 163 97 488 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=80560 $D=0
M1443 164 97 489 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=85190 $D=0
M1444 490 98 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=80560 $D=0
M1445 491 98 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=85190 $D=0
M1446 492 488 212 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=80560 $D=0
M1447 493 489 213 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=85190 $D=0
M1448 163 492 744 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=80560 $D=0
M1449 164 493 745 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=85190 $D=0
M1450 494 744 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=80560 $D=0
M1451 495 745 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=85190 $D=0
M1452 492 97 494 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=80560 $D=0
M1453 493 97 495 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=85190 $D=0
M1454 494 490 222 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=80560 $D=0
M1455 495 491 223 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=85190 $D=0
M1456 226 496 494 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=80560 $D=0
M1457 227 497 495 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=85190 $D=0
M1458 496 99 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=80560 $D=0
M1459 497 99 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=85190 $D=0
M1460 163 100 498 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=80560 $D=0
M1461 164 100 499 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=85190 $D=0
M1462 500 101 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=80560 $D=0
M1463 501 101 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=85190 $D=0
M1464 502 498 212 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=80560 $D=0
M1465 503 499 213 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=85190 $D=0
M1466 163 502 746 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=80560 $D=0
M1467 164 503 747 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=85190 $D=0
M1468 504 746 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=80560 $D=0
M1469 505 747 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=85190 $D=0
M1470 502 100 504 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=80560 $D=0
M1471 503 100 505 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=85190 $D=0
M1472 504 500 222 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=80560 $D=0
M1473 505 501 223 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=85190 $D=0
M1474 226 506 504 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=80560 $D=0
M1475 227 507 505 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=85190 $D=0
M1476 506 102 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=80560 $D=0
M1477 507 102 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=85190 $D=0
M1478 163 103 508 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=80560 $D=0
M1479 164 103 509 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=85190 $D=0
M1480 510 104 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=80560 $D=0
M1481 511 104 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=85190 $D=0
M1482 512 508 212 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=80560 $D=0
M1483 513 509 213 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=85190 $D=0
M1484 163 512 748 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=80560 $D=0
M1485 164 513 749 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=85190 $D=0
M1486 514 748 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=80560 $D=0
M1487 515 749 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=85190 $D=0
M1488 512 103 514 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=80560 $D=0
M1489 513 103 515 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=85190 $D=0
M1490 514 510 222 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=80560 $D=0
M1491 515 511 223 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=85190 $D=0
M1492 226 516 514 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=80560 $D=0
M1493 227 517 515 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=85190 $D=0
M1494 516 105 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=80560 $D=0
M1495 517 105 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=85190 $D=0
M1496 163 106 518 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=80560 $D=0
M1497 164 106 519 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=85190 $D=0
M1498 520 107 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=80560 $D=0
M1499 521 107 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=85190 $D=0
M1500 522 518 212 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=80560 $D=0
M1501 523 519 213 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=85190 $D=0
M1502 163 522 750 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=80560 $D=0
M1503 164 523 751 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=85190 $D=0
M1504 524 750 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=80560 $D=0
M1505 525 751 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=85190 $D=0
M1506 522 106 524 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=80560 $D=0
M1507 523 106 525 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=85190 $D=0
M1508 524 520 222 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=80560 $D=0
M1509 525 521 223 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=85190 $D=0
M1510 226 526 524 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=80560 $D=0
M1511 227 527 525 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=85190 $D=0
M1512 526 108 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=80560 $D=0
M1513 527 108 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=85190 $D=0
M1514 163 109 528 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=80560 $D=0
M1515 164 109 529 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=85190 $D=0
M1516 530 110 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=80560 $D=0
M1517 531 110 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=85190 $D=0
M1518 5 530 222 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=80560 $D=0
M1519 6 531 223 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=85190 $D=0
M1520 226 528 5 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=80560 $D=0
M1521 227 529 6 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=85190 $D=0
M1522 163 534 532 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=80560 $D=0
M1523 164 535 533 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=85190 $D=0
M1524 534 111 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=80560 $D=0
M1525 535 111 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=85190 $D=0
M1526 752 222 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=80560 $D=0
M1527 753 223 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=85190 $D=0
M1528 536 534 752 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=80560 $D=0
M1529 537 535 753 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=85190 $D=0
M1530 163 536 538 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=80560 $D=0
M1531 164 537 539 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=85190 $D=0
M1532 754 538 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=80560 $D=0
M1533 755 539 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=85190 $D=0
M1534 536 532 754 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=80560 $D=0
M1535 537 533 755 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=85190 $D=0
M1536 163 542 540 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=80560 $D=0
M1537 164 543 541 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=85190 $D=0
M1538 542 111 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=80560 $D=0
M1539 543 111 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=85190 $D=0
M1540 756 226 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=80560 $D=0
M1541 757 227 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=85190 $D=0
M1542 544 542 756 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=80560 $D=0
M1543 545 543 757 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=85190 $D=0
M1544 163 544 112 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=80560 $D=0
M1545 164 545 113 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=85190 $D=0
M1546 758 112 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=80560 $D=0
M1547 759 113 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=85190 $D=0
M1548 544 540 758 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=80560 $D=0
M1549 545 541 759 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=85190 $D=0
M1550 546 114 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=80560 $D=0
M1551 547 114 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=85190 $D=0
M1552 548 114 538 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=80560 $D=0
M1553 549 114 539 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=85190 $D=0
M1554 115 546 548 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=80560 $D=0
M1555 116 547 549 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=85190 $D=0
M1556 550 117 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=80560 $D=0
M1557 551 117 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=85190 $D=0
M1558 552 117 112 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=80560 $D=0
M1559 553 117 113 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=85190 $D=0
M1560 760 550 552 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=80560 $D=0
M1561 761 551 553 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=85190 $D=0
M1562 163 112 760 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=80560 $D=0
M1563 164 113 761 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=85190 $D=0
M1564 554 118 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=80560 $D=0
M1565 555 118 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=85190 $D=0
M1566 556 118 552 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=80560 $D=0
M1567 557 118 553 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=85190 $D=0
M1568 10 554 556 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=80560 $D=0
M1569 11 555 557 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=85190 $D=0
M1570 559 558 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=80560 $D=0
M1571 560 119 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=85190 $D=0
M1572 163 563 561 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=80560 $D=0
M1573 164 564 562 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=85190 $D=0
M1574 565 548 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=80560 $D=0
M1575 566 549 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=85190 $D=0
M1576 563 548 558 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=80560 $D=0
M1577 564 549 119 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=85190 $D=0
M1578 559 565 563 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=80560 $D=0
M1579 560 566 564 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=85190 $D=0
M1580 567 561 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=80560 $D=0
M1581 568 562 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=85190 $D=0
M1582 120 561 556 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=80560 $D=0
M1583 558 562 557 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=85190 $D=0
M1584 548 567 120 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=80560 $D=0
M1585 549 568 558 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=85190 $D=0
M1586 569 120 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=80560 $D=0
M1587 570 558 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=85190 $D=0
M1588 571 561 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=80560 $D=0
M1589 572 562 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=85190 $D=0
M1590 573 561 569 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=80560 $D=0
M1591 574 562 570 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=85190 $D=0
M1592 556 571 573 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=80560 $D=0
M1593 557 572 574 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=85190 $D=0
M1594 782 548 163 163 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=80200 $D=0
M1595 783 549 164 164 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=84830 $D=0
M1596 575 556 782 163 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=80200 $D=0
M1597 576 557 783 164 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=84830 $D=0
M1598 577 573 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=80560 $D=0
M1599 578 574 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=85190 $D=0
M1600 579 548 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=80560 $D=0
M1601 580 549 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=85190 $D=0
M1602 163 556 579 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=80560 $D=0
M1603 164 557 580 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=85190 $D=0
M1604 581 548 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=80560 $D=0
M1605 582 549 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=85190 $D=0
M1606 163 556 581 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=80560 $D=0
M1607 164 557 582 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=85190 $D=0
M1608 784 548 163 163 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=80380 $D=0
M1609 785 549 164 164 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=85010 $D=0
M1610 585 556 784 163 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=80380 $D=0
M1611 586 557 785 164 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=85010 $D=0
M1612 163 581 585 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=80560 $D=0
M1613 164 582 586 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=85190 $D=0
M1614 587 123 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=80560 $D=0
M1615 588 123 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=85190 $D=0
M1616 589 123 575 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=80560 $D=0
M1617 590 123 576 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=85190 $D=0
M1618 579 587 589 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=80560 $D=0
M1619 580 588 590 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=85190 $D=0
M1620 591 123 577 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=80560 $D=0
M1621 592 123 578 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=85190 $D=0
M1622 585 587 591 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=80560 $D=0
M1623 586 588 592 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=85190 $D=0
M1624 593 124 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=80560 $D=0
M1625 594 124 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=85190 $D=0
M1626 595 124 591 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=80560 $D=0
M1627 596 124 592 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=85190 $D=0
M1628 589 593 595 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=80560 $D=0
M1629 590 594 596 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=85190 $D=0
M1630 12 595 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=80560 $D=0
M1631 13 596 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=85190 $D=0
M1632 597 125 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=80560 $D=0
M1633 598 125 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=85190 $D=0
M1634 599 125 126 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=80560 $D=0
M1635 600 125 127 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=85190 $D=0
M1636 128 597 599 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=80560 $D=0
M1637 129 598 600 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=85190 $D=0
M1638 601 125 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=80560 $D=0
M1639 602 125 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=85190 $D=0
M1640 606 125 130 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=80560 $D=0
M1641 607 125 132 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=85190 $D=0
M1642 133 601 606 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=80560 $D=0
M1643 131 602 607 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=85190 $D=0
M1644 608 125 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=80560 $D=0
M1645 609 125 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=85190 $D=0
M1646 610 125 134 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=80560 $D=0
M1647 611 125 135 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=85190 $D=0
M1648 136 608 610 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=80560 $D=0
M1649 137 609 611 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=85190 $D=0
M1650 612 125 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=80560 $D=0
M1651 613 125 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=85190 $D=0
M1652 614 125 138 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=80560 $D=0
M1653 615 125 139 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=85190 $D=0
M1654 140 612 614 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=80560 $D=0
M1655 141 613 615 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=85190 $D=0
M1656 616 125 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=80560 $D=0
M1657 617 125 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=85190 $D=0
M1658 618 125 5 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=80560 $D=0
M1659 619 125 6 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=85190 $D=0
M1660 142 616 618 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=80560 $D=0
M1661 143 617 619 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=85190 $D=0
M1662 163 548 772 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=80560 $D=0
M1663 164 549 773 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=85190 $D=0
M1664 129 772 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=80560 $D=0
M1665 126 773 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=85190 $D=0
M1666 620 144 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=80560 $D=0
M1667 621 144 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=85190 $D=0
M1668 145 144 129 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=80560 $D=0
M1669 146 144 126 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=85190 $D=0
M1670 599 620 145 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=80560 $D=0
M1671 600 621 146 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=85190 $D=0
M1672 622 147 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=80560 $D=0
M1673 623 147 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=85190 $D=0
M1674 122 147 145 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=80560 $D=0
M1675 121 147 146 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=85190 $D=0
M1676 606 622 122 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=80560 $D=0
M1677 607 623 121 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=85190 $D=0
M1678 624 148 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=80560 $D=0
M1679 625 148 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=85190 $D=0
M1680 149 148 122 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=80560 $D=0
M1681 150 148 121 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=85190 $D=0
M1682 610 624 149 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=80560 $D=0
M1683 611 625 150 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=85190 $D=0
M1684 626 151 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=80560 $D=0
M1685 627 151 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=85190 $D=0
M1686 152 151 149 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=80560 $D=0
M1687 153 151 150 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=85190 $D=0
M1688 614 626 152 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=80560 $D=0
M1689 615 627 153 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=85190 $D=0
M1690 628 154 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=80560 $D=0
M1691 629 154 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=85190 $D=0
M1692 198 154 152 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=80560 $D=0
M1693 199 154 153 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=85190 $D=0
M1694 618 628 198 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=80560 $D=0
M1695 619 629 199 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=85190 $D=0
M1696 630 155 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=80560 $D=0
M1697 631 155 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=85190 $D=0
M1698 632 155 112 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=80560 $D=0
M1699 633 155 113 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=85190 $D=0
M1700 10 630 632 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=80560 $D=0
M1701 11 631 633 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=85190 $D=0
M1702 634 538 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=80560 $D=0
M1703 635 539 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=85190 $D=0
M1704 163 632 634 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=80560 $D=0
M1705 164 633 635 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=85190 $D=0
M1706 786 538 163 163 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=80380 $D=0
M1707 787 539 164 164 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=85010 $D=0
M1708 638 632 786 163 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=80380 $D=0
M1709 639 633 787 164 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=85010 $D=0
M1710 163 634 638 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=80560 $D=0
M1711 164 635 639 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=85190 $D=0
M1712 774 640 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=80560 $D=0
M1713 775 641 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=85190 $D=0
M1714 163 638 774 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=80560 $D=0
M1715 164 639 775 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=85190 $D=0
M1716 641 774 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=80560 $D=0
M1717 156 775 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=85190 $D=0
M1718 788 538 163 163 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=80200 $D=0
M1719 789 539 164 164 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=84830 $D=0
M1720 642 644 788 163 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=80200 $D=0
M1721 643 645 789 164 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=84830 $D=0
M1722 644 632 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=80560 $D=0
M1723 645 633 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=85190 $D=0
M1724 646 642 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=80560 $D=0
M1725 647 643 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=85190 $D=0
M1726 163 640 646 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=80560 $D=0
M1727 164 641 647 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=85190 $D=0
M1728 649 157 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=80560 $D=0
M1729 650 648 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=85190 $D=0
M1730 648 646 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=80560 $D=0
M1731 158 647 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=85190 $D=0
M1732 163 649 648 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=80560 $D=0
M1733 164 650 158 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=85190 $D=0
M1734 652 651 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=80560 $D=0
M1735 653 159 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=85190 $D=0
M1736 163 656 654 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=80560 $D=0
M1737 164 657 655 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=85190 $D=0
M1738 658 115 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=80560 $D=0
M1739 659 116 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=85190 $D=0
M1740 656 115 651 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=80560 $D=0
M1741 657 116 159 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=85190 $D=0
M1742 652 658 656 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=80560 $D=0
M1743 653 659 657 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=85190 $D=0
M1744 660 654 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=80560 $D=0
M1745 661 655 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=85190 $D=0
M1746 160 654 5 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=80560 $D=0
M1747 651 655 6 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=85190 $D=0
M1748 115 660 160 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=80560 $D=0
M1749 116 661 651 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=85190 $D=0
M1750 662 160 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=80560 $D=0
M1751 663 651 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=85190 $D=0
M1752 664 654 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=80560 $D=0
M1753 665 655 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=85190 $D=0
M1754 200 654 662 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=80560 $D=0
M1755 201 655 663 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=85190 $D=0
M1756 5 664 200 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=80560 $D=0
M1757 6 665 201 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=85190 $D=0
M1758 666 161 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=80560 $D=0
M1759 667 161 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=85190 $D=0
M1760 668 161 200 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=80560 $D=0
M1761 669 161 201 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=85190 $D=0
M1762 12 666 668 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=80560 $D=0
M1763 13 667 669 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=85190 $D=0
M1764 670 162 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=80560 $D=0
M1765 671 162 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=85190 $D=0
M1766 162 162 668 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=80560 $D=0
M1767 162 162 669 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=85190 $D=0
M1768 5 670 162 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=80560 $D=0
M1769 6 671 162 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=85190 $D=0
M1770 672 111 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=80560 $D=0
M1771 673 111 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=85190 $D=0
M1772 163 672 674 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=80560 $D=0
M1773 164 673 675 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=85190 $D=0
M1774 676 111 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=80560 $D=0
M1775 677 111 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=85190 $D=0
M1776 678 674 162 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=80560 $D=0
M1777 679 675 162 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=85190 $D=0
M1778 163 678 776 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=80560 $D=0
M1779 164 679 777 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=85190 $D=0
M1780 680 776 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=80560 $D=0
M1781 681 777 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=85190 $D=0
M1782 678 672 680 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=80560 $D=0
M1783 679 673 681 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=85190 $D=0
M1784 682 676 680 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=80560 $D=0
M1785 683 677 681 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=85190 $D=0
M1786 163 686 684 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=80560 $D=0
M1787 164 687 685 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=85190 $D=0
M1788 686 111 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=80560 $D=0
M1789 687 111 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=85190 $D=0
M1790 778 682 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=80560 $D=0
M1791 779 683 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=85190 $D=0
M1792 688 686 778 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=80560 $D=0
M1793 689 687 779 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=85190 $D=0
M1794 163 688 115 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=80560 $D=0
M1795 164 689 116 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=85190 $D=0
M1796 780 115 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=80560 $D=0
M1797 781 116 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=85190 $D=0
M1798 688 684 780 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=80560 $D=0
M1799 689 685 781 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=85190 $D=0
.ENDS
***************************************
.SUBCKT ICV_31 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141
+ 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161
+ 162 163 164 165 166
** N=799 EP=165 IP=1514 FDC=1800
M0 176 1 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=70050 $D=1
M1 177 1 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=74680 $D=1
M2 178 176 2 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=70050 $D=1
M3 179 177 3 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=74680 $D=1
M4 5 1 178 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=70050 $D=1
M5 6 1 179 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=74680 $D=1
M6 180 176 4 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=70050 $D=1
M7 181 177 4 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=74680 $D=1
M8 3 1 180 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=70050 $D=1
M9 3 1 181 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=74680 $D=1
M10 182 176 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=70050 $D=1
M11 183 177 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=74680 $D=1
M12 5 1 182 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=70050 $D=1
M13 3 1 183 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=74680 $D=1
M14 186 184 182 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=70050 $D=1
M15 187 185 183 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=74680 $D=1
M16 184 7 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=70050 $D=1
M17 185 7 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=74680 $D=1
M18 188 184 180 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=70050 $D=1
M19 189 185 181 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=74680 $D=1
M20 178 7 188 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=70050 $D=1
M21 179 7 189 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=74680 $D=1
M22 190 8 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=70050 $D=1
M23 191 8 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=74680 $D=1
M24 192 190 188 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=70050 $D=1
M25 193 191 189 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=74680 $D=1
M26 186 8 192 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=70050 $D=1
M27 187 8 193 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=74680 $D=1
M28 194 9 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=70050 $D=1
M29 195 9 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=74680 $D=1
M30 196 194 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=70050 $D=1
M31 197 195 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=74680 $D=1
M32 10 9 196 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=70050 $D=1
M33 11 9 197 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=74680 $D=1
M34 198 194 12 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=70050 $D=1
M35 199 195 13 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=74680 $D=1
M36 14 9 198 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=70050 $D=1
M37 200 9 199 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=74680 $D=1
M38 203 194 201 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=70050 $D=1
M39 204 195 202 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=74680 $D=1
M40 192 9 203 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=70050 $D=1
M41 193 9 204 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=74680 $D=1
M42 207 205 203 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=70050 $D=1
M43 208 206 204 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=74680 $D=1
M44 205 15 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=70050 $D=1
M45 206 15 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=74680 $D=1
M46 209 205 198 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=70050 $D=1
M47 210 206 199 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=74680 $D=1
M48 196 15 209 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=70050 $D=1
M49 197 15 210 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=74680 $D=1
M50 211 16 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=70050 $D=1
M51 212 16 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=74680 $D=1
M52 213 211 209 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=70050 $D=1
M53 214 212 210 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=74680 $D=1
M54 207 16 213 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=70050 $D=1
M55 208 16 214 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=74680 $D=1
M56 5 17 215 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=70050 $D=1
M57 6 17 216 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=74680 $D=1
M58 217 18 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=70050 $D=1
M59 218 18 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=74680 $D=1
M60 219 17 213 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=70050 $D=1
M61 220 17 214 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=74680 $D=1
M62 5 219 690 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=70050 $D=1
M63 6 220 691 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=74680 $D=1
M64 221 690 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=70050 $D=1
M65 222 691 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=74680 $D=1
M66 219 215 221 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=70050 $D=1
M67 220 216 222 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=74680 $D=1
M68 221 18 223 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=70050 $D=1
M69 222 18 224 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=74680 $D=1
M70 227 19 221 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=70050 $D=1
M71 228 19 222 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=74680 $D=1
M72 225 19 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=70050 $D=1
M73 226 19 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=74680 $D=1
M74 5 20 229 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=70050 $D=1
M75 6 20 230 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=74680 $D=1
M76 231 21 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=70050 $D=1
M77 232 21 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=74680 $D=1
M78 233 20 213 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=70050 $D=1
M79 234 20 214 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=74680 $D=1
M80 5 233 692 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=70050 $D=1
M81 6 234 693 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=74680 $D=1
M82 235 692 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=70050 $D=1
M83 236 693 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=74680 $D=1
M84 233 229 235 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=70050 $D=1
M85 234 230 236 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=74680 $D=1
M86 235 21 223 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=70050 $D=1
M87 236 21 224 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=74680 $D=1
M88 227 22 235 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=70050 $D=1
M89 228 22 236 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=74680 $D=1
M90 237 22 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=70050 $D=1
M91 238 22 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=74680 $D=1
M92 5 23 239 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=70050 $D=1
M93 6 23 240 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=74680 $D=1
M94 241 24 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=70050 $D=1
M95 242 24 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=74680 $D=1
M96 243 23 213 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=70050 $D=1
M97 244 23 214 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=74680 $D=1
M98 5 243 694 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=70050 $D=1
M99 6 244 695 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=74680 $D=1
M100 245 694 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=70050 $D=1
M101 246 695 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=74680 $D=1
M102 243 239 245 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=70050 $D=1
M103 244 240 246 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=74680 $D=1
M104 245 24 223 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=70050 $D=1
M105 246 24 224 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=74680 $D=1
M106 227 25 245 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=70050 $D=1
M107 228 25 246 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=74680 $D=1
M108 247 25 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=70050 $D=1
M109 248 25 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=74680 $D=1
M110 5 26 249 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=70050 $D=1
M111 6 26 250 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=74680 $D=1
M112 251 27 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=70050 $D=1
M113 252 27 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=74680 $D=1
M114 253 26 213 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=70050 $D=1
M115 254 26 214 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=74680 $D=1
M116 5 253 696 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=70050 $D=1
M117 6 254 697 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=74680 $D=1
M118 255 696 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=70050 $D=1
M119 256 697 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=74680 $D=1
M120 253 249 255 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=70050 $D=1
M121 254 250 256 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=74680 $D=1
M122 255 27 223 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=70050 $D=1
M123 256 27 224 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=74680 $D=1
M124 227 28 255 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=70050 $D=1
M125 228 28 256 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=74680 $D=1
M126 257 28 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=70050 $D=1
M127 258 28 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=74680 $D=1
M128 5 29 259 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=70050 $D=1
M129 6 29 260 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=74680 $D=1
M130 261 30 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=70050 $D=1
M131 262 30 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=74680 $D=1
M132 263 29 213 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=70050 $D=1
M133 264 29 214 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=74680 $D=1
M134 5 263 698 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=70050 $D=1
M135 6 264 699 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=74680 $D=1
M136 265 698 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=70050 $D=1
M137 266 699 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=74680 $D=1
M138 263 259 265 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=70050 $D=1
M139 264 260 266 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=74680 $D=1
M140 265 30 223 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=70050 $D=1
M141 266 30 224 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=74680 $D=1
M142 227 31 265 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=70050 $D=1
M143 228 31 266 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=74680 $D=1
M144 267 31 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=70050 $D=1
M145 268 31 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=74680 $D=1
M146 5 32 269 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=70050 $D=1
M147 6 32 270 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=74680 $D=1
M148 271 33 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=70050 $D=1
M149 272 33 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=74680 $D=1
M150 273 32 213 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=70050 $D=1
M151 274 32 214 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=74680 $D=1
M152 5 273 700 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=70050 $D=1
M153 6 274 701 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=74680 $D=1
M154 275 700 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=70050 $D=1
M155 276 701 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=74680 $D=1
M156 273 269 275 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=70050 $D=1
M157 274 270 276 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=74680 $D=1
M158 275 33 223 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=70050 $D=1
M159 276 33 224 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=74680 $D=1
M160 227 34 275 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=70050 $D=1
M161 228 34 276 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=74680 $D=1
M162 277 34 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=70050 $D=1
M163 278 34 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=74680 $D=1
M164 5 35 279 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=70050 $D=1
M165 6 35 280 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=74680 $D=1
M166 281 36 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=70050 $D=1
M167 282 36 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=74680 $D=1
M168 283 35 213 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=70050 $D=1
M169 284 35 214 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=74680 $D=1
M170 5 283 702 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=70050 $D=1
M171 6 284 703 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=74680 $D=1
M172 285 702 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=70050 $D=1
M173 286 703 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=74680 $D=1
M174 283 279 285 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=70050 $D=1
M175 284 280 286 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=74680 $D=1
M176 285 36 223 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=70050 $D=1
M177 286 36 224 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=74680 $D=1
M178 227 37 285 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=70050 $D=1
M179 228 37 286 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=74680 $D=1
M180 287 37 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=70050 $D=1
M181 288 37 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=74680 $D=1
M182 5 38 289 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=70050 $D=1
M183 6 38 290 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=74680 $D=1
M184 291 39 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=70050 $D=1
M185 292 39 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=74680 $D=1
M186 293 38 213 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=70050 $D=1
M187 294 38 214 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=74680 $D=1
M188 5 293 704 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=70050 $D=1
M189 6 294 705 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=74680 $D=1
M190 295 704 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=70050 $D=1
M191 296 705 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=74680 $D=1
M192 293 289 295 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=70050 $D=1
M193 294 290 296 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=74680 $D=1
M194 295 39 223 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=70050 $D=1
M195 296 39 224 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=74680 $D=1
M196 227 40 295 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=70050 $D=1
M197 228 40 296 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=74680 $D=1
M198 297 40 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=70050 $D=1
M199 298 40 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=74680 $D=1
M200 5 41 299 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=70050 $D=1
M201 6 41 300 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=74680 $D=1
M202 301 42 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=70050 $D=1
M203 302 42 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=74680 $D=1
M204 303 41 213 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=70050 $D=1
M205 304 41 214 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=74680 $D=1
M206 5 303 706 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=70050 $D=1
M207 6 304 707 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=74680 $D=1
M208 305 706 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=70050 $D=1
M209 306 707 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=74680 $D=1
M210 303 299 305 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=70050 $D=1
M211 304 300 306 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=74680 $D=1
M212 305 42 223 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=70050 $D=1
M213 306 42 224 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=74680 $D=1
M214 227 43 305 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=70050 $D=1
M215 228 43 306 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=74680 $D=1
M216 307 43 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=70050 $D=1
M217 308 43 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=74680 $D=1
M218 5 44 309 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=70050 $D=1
M219 6 44 310 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=74680 $D=1
M220 311 45 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=70050 $D=1
M221 312 45 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=74680 $D=1
M222 313 44 213 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=70050 $D=1
M223 314 44 214 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=74680 $D=1
M224 5 313 708 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=70050 $D=1
M225 6 314 709 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=74680 $D=1
M226 315 708 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=70050 $D=1
M227 316 709 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=74680 $D=1
M228 313 309 315 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=70050 $D=1
M229 314 310 316 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=74680 $D=1
M230 315 45 223 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=70050 $D=1
M231 316 45 224 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=74680 $D=1
M232 227 46 315 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=70050 $D=1
M233 228 46 316 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=74680 $D=1
M234 317 46 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=70050 $D=1
M235 318 46 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=74680 $D=1
M236 5 47 319 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=70050 $D=1
M237 6 47 320 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=74680 $D=1
M238 321 48 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=70050 $D=1
M239 322 48 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=74680 $D=1
M240 323 47 213 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=70050 $D=1
M241 324 47 214 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=74680 $D=1
M242 5 323 710 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=70050 $D=1
M243 6 324 711 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=74680 $D=1
M244 325 710 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=70050 $D=1
M245 326 711 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=74680 $D=1
M246 323 319 325 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=70050 $D=1
M247 324 320 326 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=74680 $D=1
M248 325 48 223 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=70050 $D=1
M249 326 48 224 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=74680 $D=1
M250 227 49 325 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=70050 $D=1
M251 228 49 326 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=74680 $D=1
M252 327 49 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=70050 $D=1
M253 328 49 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=74680 $D=1
M254 5 50 329 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=70050 $D=1
M255 6 50 330 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=74680 $D=1
M256 331 51 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=70050 $D=1
M257 332 51 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=74680 $D=1
M258 333 50 213 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=70050 $D=1
M259 334 50 214 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=74680 $D=1
M260 5 333 712 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=70050 $D=1
M261 6 334 713 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=74680 $D=1
M262 335 712 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=70050 $D=1
M263 336 713 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=74680 $D=1
M264 333 329 335 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=70050 $D=1
M265 334 330 336 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=74680 $D=1
M266 335 51 223 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=70050 $D=1
M267 336 51 224 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=74680 $D=1
M268 227 52 335 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=70050 $D=1
M269 228 52 336 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=74680 $D=1
M270 337 52 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=70050 $D=1
M271 338 52 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=74680 $D=1
M272 5 53 339 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=70050 $D=1
M273 6 53 340 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=74680 $D=1
M274 341 54 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=70050 $D=1
M275 342 54 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=74680 $D=1
M276 343 53 213 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=70050 $D=1
M277 344 53 214 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=74680 $D=1
M278 5 343 714 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=70050 $D=1
M279 6 344 715 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=74680 $D=1
M280 345 714 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=70050 $D=1
M281 346 715 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=74680 $D=1
M282 343 339 345 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=70050 $D=1
M283 344 340 346 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=74680 $D=1
M284 345 54 223 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=70050 $D=1
M285 346 54 224 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=74680 $D=1
M286 227 55 345 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=70050 $D=1
M287 228 55 346 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=74680 $D=1
M288 347 55 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=70050 $D=1
M289 348 55 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=74680 $D=1
M290 5 56 349 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=70050 $D=1
M291 6 56 350 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=74680 $D=1
M292 351 57 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=70050 $D=1
M293 352 57 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=74680 $D=1
M294 353 56 213 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=70050 $D=1
M295 354 56 214 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=74680 $D=1
M296 5 353 716 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=70050 $D=1
M297 6 354 717 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=74680 $D=1
M298 355 716 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=70050 $D=1
M299 356 717 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=74680 $D=1
M300 353 349 355 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=70050 $D=1
M301 354 350 356 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=74680 $D=1
M302 355 57 223 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=70050 $D=1
M303 356 57 224 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=74680 $D=1
M304 227 58 355 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=70050 $D=1
M305 228 58 356 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=74680 $D=1
M306 357 58 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=70050 $D=1
M307 358 58 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=74680 $D=1
M308 5 59 359 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=70050 $D=1
M309 6 59 360 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=74680 $D=1
M310 361 60 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=70050 $D=1
M311 362 60 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=74680 $D=1
M312 363 59 213 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=70050 $D=1
M313 364 59 214 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=74680 $D=1
M314 5 363 718 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=70050 $D=1
M315 6 364 719 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=74680 $D=1
M316 365 718 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=70050 $D=1
M317 366 719 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=74680 $D=1
M318 363 359 365 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=70050 $D=1
M319 364 360 366 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=74680 $D=1
M320 365 60 223 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=70050 $D=1
M321 366 60 224 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=74680 $D=1
M322 227 61 365 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=70050 $D=1
M323 228 61 366 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=74680 $D=1
M324 367 61 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=70050 $D=1
M325 368 61 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=74680 $D=1
M326 5 62 369 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=70050 $D=1
M327 6 62 370 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=74680 $D=1
M328 371 63 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=70050 $D=1
M329 372 63 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=74680 $D=1
M330 373 62 213 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=70050 $D=1
M331 374 62 214 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=74680 $D=1
M332 5 373 720 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=70050 $D=1
M333 6 374 721 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=74680 $D=1
M334 375 720 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=70050 $D=1
M335 376 721 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=74680 $D=1
M336 373 369 375 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=70050 $D=1
M337 374 370 376 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=74680 $D=1
M338 375 63 223 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=70050 $D=1
M339 376 63 224 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=74680 $D=1
M340 227 64 375 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=70050 $D=1
M341 228 64 376 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=74680 $D=1
M342 377 64 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=70050 $D=1
M343 378 64 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=74680 $D=1
M344 5 65 379 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=70050 $D=1
M345 6 65 380 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=74680 $D=1
M346 381 66 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=70050 $D=1
M347 382 66 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=74680 $D=1
M348 383 65 213 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=70050 $D=1
M349 384 65 214 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=74680 $D=1
M350 5 383 722 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=70050 $D=1
M351 6 384 723 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=74680 $D=1
M352 385 722 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=70050 $D=1
M353 386 723 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=74680 $D=1
M354 383 379 385 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=70050 $D=1
M355 384 380 386 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=74680 $D=1
M356 385 66 223 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=70050 $D=1
M357 386 66 224 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=74680 $D=1
M358 227 67 385 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=70050 $D=1
M359 228 67 386 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=74680 $D=1
M360 387 67 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=70050 $D=1
M361 388 67 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=74680 $D=1
M362 5 68 389 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=70050 $D=1
M363 6 68 390 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=74680 $D=1
M364 391 69 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=70050 $D=1
M365 392 69 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=74680 $D=1
M366 393 68 213 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=70050 $D=1
M367 394 68 214 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=74680 $D=1
M368 5 393 724 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=70050 $D=1
M369 6 394 725 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=74680 $D=1
M370 395 724 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=70050 $D=1
M371 396 725 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=74680 $D=1
M372 393 389 395 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=70050 $D=1
M373 394 390 396 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=74680 $D=1
M374 395 69 223 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=70050 $D=1
M375 396 69 224 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=74680 $D=1
M376 227 70 395 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=70050 $D=1
M377 228 70 396 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=74680 $D=1
M378 397 70 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=70050 $D=1
M379 398 70 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=74680 $D=1
M380 5 71 399 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=70050 $D=1
M381 6 71 400 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=74680 $D=1
M382 401 72 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=70050 $D=1
M383 402 72 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=74680 $D=1
M384 403 71 213 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=70050 $D=1
M385 404 71 214 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=74680 $D=1
M386 5 403 726 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=70050 $D=1
M387 6 404 727 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=74680 $D=1
M388 405 726 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=70050 $D=1
M389 406 727 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=74680 $D=1
M390 403 399 405 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=70050 $D=1
M391 404 400 406 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=74680 $D=1
M392 405 72 223 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=70050 $D=1
M393 406 72 224 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=74680 $D=1
M394 227 73 405 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=70050 $D=1
M395 228 73 406 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=74680 $D=1
M396 407 73 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=70050 $D=1
M397 408 73 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=74680 $D=1
M398 5 74 409 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=70050 $D=1
M399 6 74 410 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=74680 $D=1
M400 411 75 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=70050 $D=1
M401 412 75 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=74680 $D=1
M402 413 74 213 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=70050 $D=1
M403 414 74 214 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=74680 $D=1
M404 5 413 728 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=70050 $D=1
M405 6 414 729 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=74680 $D=1
M406 415 728 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=70050 $D=1
M407 416 729 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=74680 $D=1
M408 413 409 415 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=70050 $D=1
M409 414 410 416 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=74680 $D=1
M410 415 75 223 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=70050 $D=1
M411 416 75 224 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=74680 $D=1
M412 227 76 415 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=70050 $D=1
M413 228 76 416 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=74680 $D=1
M414 417 76 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=70050 $D=1
M415 418 76 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=74680 $D=1
M416 5 77 419 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=70050 $D=1
M417 6 77 420 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=74680 $D=1
M418 421 78 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=70050 $D=1
M419 422 78 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=74680 $D=1
M420 423 77 213 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=70050 $D=1
M421 424 77 214 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=74680 $D=1
M422 5 423 730 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=70050 $D=1
M423 6 424 731 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=74680 $D=1
M424 425 730 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=70050 $D=1
M425 426 731 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=74680 $D=1
M426 423 419 425 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=70050 $D=1
M427 424 420 426 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=74680 $D=1
M428 425 78 223 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=70050 $D=1
M429 426 78 224 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=74680 $D=1
M430 227 79 425 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=70050 $D=1
M431 228 79 426 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=74680 $D=1
M432 427 79 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=70050 $D=1
M433 428 79 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=74680 $D=1
M434 5 80 429 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=70050 $D=1
M435 6 80 430 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=74680 $D=1
M436 431 81 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=70050 $D=1
M437 432 81 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=74680 $D=1
M438 433 80 213 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=70050 $D=1
M439 434 80 214 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=74680 $D=1
M440 5 433 732 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=70050 $D=1
M441 6 434 733 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=74680 $D=1
M442 435 732 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=70050 $D=1
M443 436 733 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=74680 $D=1
M444 433 429 435 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=70050 $D=1
M445 434 430 436 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=74680 $D=1
M446 435 81 223 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=70050 $D=1
M447 436 81 224 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=74680 $D=1
M448 227 82 435 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=70050 $D=1
M449 228 82 436 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=74680 $D=1
M450 437 82 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=70050 $D=1
M451 438 82 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=74680 $D=1
M452 5 83 439 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=70050 $D=1
M453 6 83 440 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=74680 $D=1
M454 441 84 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=70050 $D=1
M455 442 84 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=74680 $D=1
M456 443 83 213 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=70050 $D=1
M457 444 83 214 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=74680 $D=1
M458 5 443 734 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=70050 $D=1
M459 6 444 735 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=74680 $D=1
M460 445 734 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=70050 $D=1
M461 446 735 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=74680 $D=1
M462 443 439 445 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=70050 $D=1
M463 444 440 446 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=74680 $D=1
M464 445 84 223 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=70050 $D=1
M465 446 84 224 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=74680 $D=1
M466 227 85 445 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=70050 $D=1
M467 228 85 446 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=74680 $D=1
M468 447 85 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=70050 $D=1
M469 448 85 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=74680 $D=1
M470 5 86 449 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=70050 $D=1
M471 6 86 450 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=74680 $D=1
M472 451 87 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=70050 $D=1
M473 452 87 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=74680 $D=1
M474 453 86 213 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=70050 $D=1
M475 454 86 214 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=74680 $D=1
M476 5 453 736 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=70050 $D=1
M477 6 454 737 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=74680 $D=1
M478 455 736 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=70050 $D=1
M479 456 737 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=74680 $D=1
M480 453 449 455 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=70050 $D=1
M481 454 450 456 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=74680 $D=1
M482 455 87 223 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=70050 $D=1
M483 456 87 224 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=74680 $D=1
M484 227 88 455 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=70050 $D=1
M485 228 88 456 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=74680 $D=1
M486 457 88 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=70050 $D=1
M487 458 88 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=74680 $D=1
M488 5 89 459 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=70050 $D=1
M489 6 89 460 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=74680 $D=1
M490 461 90 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=70050 $D=1
M491 462 90 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=74680 $D=1
M492 463 89 213 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=70050 $D=1
M493 464 89 214 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=74680 $D=1
M494 5 463 738 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=70050 $D=1
M495 6 464 739 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=74680 $D=1
M496 465 738 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=70050 $D=1
M497 466 739 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=74680 $D=1
M498 463 459 465 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=70050 $D=1
M499 464 460 466 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=74680 $D=1
M500 465 90 223 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=70050 $D=1
M501 466 90 224 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=74680 $D=1
M502 227 91 465 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=70050 $D=1
M503 228 91 466 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=74680 $D=1
M504 467 91 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=70050 $D=1
M505 468 91 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=74680 $D=1
M506 5 92 469 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=70050 $D=1
M507 6 92 470 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=74680 $D=1
M508 471 93 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=70050 $D=1
M509 472 93 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=74680 $D=1
M510 473 92 213 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=70050 $D=1
M511 474 92 214 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=74680 $D=1
M512 5 473 740 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=70050 $D=1
M513 6 474 741 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=74680 $D=1
M514 475 740 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=70050 $D=1
M515 476 741 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=74680 $D=1
M516 473 469 475 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=70050 $D=1
M517 474 470 476 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=74680 $D=1
M518 475 93 223 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=70050 $D=1
M519 476 93 224 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=74680 $D=1
M520 227 94 475 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=70050 $D=1
M521 228 94 476 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=74680 $D=1
M522 477 94 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=70050 $D=1
M523 478 94 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=74680 $D=1
M524 5 95 479 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=70050 $D=1
M525 6 95 480 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=74680 $D=1
M526 481 96 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=70050 $D=1
M527 482 96 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=74680 $D=1
M528 483 95 213 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=70050 $D=1
M529 484 95 214 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=74680 $D=1
M530 5 483 742 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=70050 $D=1
M531 6 484 743 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=74680 $D=1
M532 485 742 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=70050 $D=1
M533 486 743 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=74680 $D=1
M534 483 479 485 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=70050 $D=1
M535 484 480 486 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=74680 $D=1
M536 485 96 223 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=70050 $D=1
M537 486 96 224 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=74680 $D=1
M538 227 97 485 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=70050 $D=1
M539 228 97 486 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=74680 $D=1
M540 487 97 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=70050 $D=1
M541 488 97 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=74680 $D=1
M542 5 98 489 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=70050 $D=1
M543 6 98 490 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=74680 $D=1
M544 491 99 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=70050 $D=1
M545 492 99 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=74680 $D=1
M546 493 98 213 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=70050 $D=1
M547 494 98 214 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=74680 $D=1
M548 5 493 744 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=70050 $D=1
M549 6 494 745 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=74680 $D=1
M550 495 744 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=70050 $D=1
M551 496 745 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=74680 $D=1
M552 493 489 495 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=70050 $D=1
M553 494 490 496 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=74680 $D=1
M554 495 99 223 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=70050 $D=1
M555 496 99 224 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=74680 $D=1
M556 227 100 495 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=70050 $D=1
M557 228 100 496 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=74680 $D=1
M558 497 100 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=70050 $D=1
M559 498 100 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=74680 $D=1
M560 5 101 499 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=70050 $D=1
M561 6 101 500 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=74680 $D=1
M562 501 102 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=70050 $D=1
M563 502 102 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=74680 $D=1
M564 503 101 213 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=70050 $D=1
M565 504 101 214 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=74680 $D=1
M566 5 503 746 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=70050 $D=1
M567 6 504 747 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=74680 $D=1
M568 505 746 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=70050 $D=1
M569 506 747 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=74680 $D=1
M570 503 499 505 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=70050 $D=1
M571 504 500 506 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=74680 $D=1
M572 505 102 223 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=70050 $D=1
M573 506 102 224 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=74680 $D=1
M574 227 103 505 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=70050 $D=1
M575 228 103 506 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=74680 $D=1
M576 507 103 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=70050 $D=1
M577 508 103 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=74680 $D=1
M578 5 104 509 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=70050 $D=1
M579 6 104 510 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=74680 $D=1
M580 511 105 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=70050 $D=1
M581 512 105 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=74680 $D=1
M582 513 104 213 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=70050 $D=1
M583 514 104 214 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=74680 $D=1
M584 5 513 748 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=70050 $D=1
M585 6 514 749 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=74680 $D=1
M586 515 748 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=70050 $D=1
M587 516 749 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=74680 $D=1
M588 513 509 515 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=70050 $D=1
M589 514 510 516 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=74680 $D=1
M590 515 105 223 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=70050 $D=1
M591 516 105 224 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=74680 $D=1
M592 227 106 515 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=70050 $D=1
M593 228 106 516 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=74680 $D=1
M594 517 106 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=70050 $D=1
M595 518 106 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=74680 $D=1
M596 5 107 519 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=70050 $D=1
M597 6 107 520 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=74680 $D=1
M598 521 108 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=70050 $D=1
M599 522 108 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=74680 $D=1
M600 523 107 213 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=70050 $D=1
M601 524 107 214 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=74680 $D=1
M602 5 523 750 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=70050 $D=1
M603 6 524 751 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=74680 $D=1
M604 525 750 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=70050 $D=1
M605 526 751 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=74680 $D=1
M606 523 519 525 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=70050 $D=1
M607 524 520 526 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=74680 $D=1
M608 525 108 223 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=70050 $D=1
M609 526 108 224 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=74680 $D=1
M610 227 109 525 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=70050 $D=1
M611 228 109 526 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=74680 $D=1
M612 527 109 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=70050 $D=1
M613 528 109 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=74680 $D=1
M614 5 110 529 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=70050 $D=1
M615 6 110 530 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=74680 $D=1
M616 531 111 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=70050 $D=1
M617 532 111 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=74680 $D=1
M618 5 111 223 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=70050 $D=1
M619 6 111 224 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=74680 $D=1
M620 227 110 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=70050 $D=1
M621 228 110 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=74680 $D=1
M622 5 535 533 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=70050 $D=1
M623 6 536 534 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=74680 $D=1
M624 535 112 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=70050 $D=1
M625 536 112 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=74680 $D=1
M626 752 223 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=70050 $D=1
M627 753 224 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=74680 $D=1
M628 537 533 752 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=70050 $D=1
M629 538 534 753 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=74680 $D=1
M630 5 537 539 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=70050 $D=1
M631 6 538 540 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=74680 $D=1
M632 754 539 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=70050 $D=1
M633 755 540 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=74680 $D=1
M634 537 535 754 5 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=70050 $D=1
M635 538 536 755 6 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=74680 $D=1
M636 5 543 541 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=70050 $D=1
M637 6 544 542 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=74680 $D=1
M638 543 112 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=70050 $D=1
M639 544 112 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=74680 $D=1
M640 756 227 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=70050 $D=1
M641 757 228 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=74680 $D=1
M642 545 541 756 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=70050 $D=1
M643 546 542 757 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=74680 $D=1
M644 5 545 113 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=70050 $D=1
M645 6 546 114 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=74680 $D=1
M646 758 113 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=70050 $D=1
M647 759 114 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=74680 $D=1
M648 545 543 758 5 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=70050 $D=1
M649 546 544 759 6 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=74680 $D=1
M650 547 115 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=70050 $D=1
M651 548 115 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=74680 $D=1
M652 549 547 539 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=70050 $D=1
M653 550 548 540 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=74680 $D=1
M654 116 115 549 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=70050 $D=1
M655 117 115 550 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=74680 $D=1
M656 551 118 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=70050 $D=1
M657 552 118 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=74680 $D=1
M658 553 551 113 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=70050 $D=1
M659 554 552 114 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=74680 $D=1
M660 760 118 553 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=70050 $D=1
M661 761 118 554 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=74680 $D=1
M662 5 113 760 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=70050 $D=1
M663 6 114 761 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=74680 $D=1
M664 555 119 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=70050 $D=1
M665 556 119 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=74680 $D=1
M666 557 555 553 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=70050 $D=1
M667 558 556 554 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=74680 $D=1
M668 10 119 557 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=70050 $D=1
M669 11 119 558 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=74680 $D=1
M670 560 559 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=70050 $D=1
M671 561 120 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=74680 $D=1
M672 5 564 562 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=70050 $D=1
M673 6 565 563 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=74680 $D=1
M674 566 549 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=70050 $D=1
M675 567 550 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=74680 $D=1
M676 564 566 559 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=70050 $D=1
M677 565 567 120 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=74680 $D=1
M678 560 549 564 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=70050 $D=1
M679 561 550 565 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=74680 $D=1
M680 568 562 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=70050 $D=1
M681 569 563 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=74680 $D=1
M682 570 568 557 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=70050 $D=1
M683 559 569 558 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=74680 $D=1
M684 549 562 570 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=70050 $D=1
M685 550 563 559 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=74680 $D=1
M686 571 570 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=70050 $D=1
M687 572 559 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=74680 $D=1
M688 573 562 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=70050 $D=1
M689 574 563 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=74680 $D=1
M690 575 573 571 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=70050 $D=1
M691 576 574 572 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=74680 $D=1
M692 557 562 575 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=70050 $D=1
M693 558 563 576 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=74680 $D=1
M694 577 549 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=70050 $D=1
M695 578 550 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=74680 $D=1
M696 5 557 577 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=70050 $D=1
M697 6 558 578 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=74680 $D=1
M698 579 575 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=70050 $D=1
M699 580 576 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=74680 $D=1
M700 788 549 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=70050 $D=1
M701 789 550 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=74680 $D=1
M702 581 557 788 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=70050 $D=1
M703 582 558 789 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=74680 $D=1
M704 790 549 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=70050 $D=1
M705 791 550 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=74680 $D=1
M706 583 557 790 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=70050 $D=1
M707 584 558 791 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=74680 $D=1
M708 587 549 585 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=70050 $D=1
M709 588 550 586 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=74680 $D=1
M710 585 557 587 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=70050 $D=1
M711 586 558 588 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=74680 $D=1
M712 5 583 585 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=70050 $D=1
M713 6 584 586 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=74680 $D=1
M714 589 125 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=70050 $D=1
M715 590 125 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=74680 $D=1
M716 591 589 577 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=70050 $D=1
M717 592 590 578 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=74680 $D=1
M718 581 125 591 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=70050 $D=1
M719 582 125 592 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=74680 $D=1
M720 593 589 579 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=70050 $D=1
M721 594 590 580 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=74680 $D=1
M722 587 125 593 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=70050 $D=1
M723 588 125 594 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=74680 $D=1
M724 595 126 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=70050 $D=1
M725 596 126 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=74680 $D=1
M726 597 595 593 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=70050 $D=1
M727 598 596 594 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=74680 $D=1
M728 591 126 597 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=70050 $D=1
M729 592 126 598 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=74680 $D=1
M730 12 597 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=70050 $D=1
M731 13 598 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=74680 $D=1
M732 599 127 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=70050 $D=1
M733 600 127 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=74680 $D=1
M734 601 599 128 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=70050 $D=1
M735 602 600 129 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=74680 $D=1
M736 130 127 601 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=70050 $D=1
M737 131 127 602 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=74680 $D=1
M738 603 127 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=70050 $D=1
M739 604 127 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=74680 $D=1
M740 606 603 132 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=70050 $D=1
M741 607 604 133 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=74680 $D=1
M742 134 127 606 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=70050 $D=1
M743 135 127 607 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=74680 $D=1
M744 608 127 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=70050 $D=1
M745 609 127 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=74680 $D=1
M746 610 608 122 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=70050 $D=1
M747 611 609 136 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=74680 $D=1
M748 137 127 610 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=70050 $D=1
M749 138 127 611 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=74680 $D=1
M750 612 127 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=70050 $D=1
M751 613 127 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=74680 $D=1
M752 614 612 139 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=70050 $D=1
M753 615 613 140 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=74680 $D=1
M754 141 127 614 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=70050 $D=1
M755 142 127 615 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=74680 $D=1
M756 616 127 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=70050 $D=1
M757 617 127 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=74680 $D=1
M758 618 616 143 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=70050 $D=1
M759 619 617 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=74680 $D=1
M760 144 127 618 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=70050 $D=1
M761 145 127 619 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=74680 $D=1
M762 5 549 770 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=70050 $D=1
M763 6 550 771 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=74680 $D=1
M764 131 770 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=70050 $D=1
M765 128 771 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=74680 $D=1
M766 620 146 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=70050 $D=1
M767 621 146 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=74680 $D=1
M768 147 620 131 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=70050 $D=1
M769 148 621 128 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=74680 $D=1
M770 601 146 147 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=70050 $D=1
M771 602 146 148 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=74680 $D=1
M772 622 149 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=70050 $D=1
M773 623 149 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=74680 $D=1
M774 121 622 147 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=70050 $D=1
M775 124 623 148 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=74680 $D=1
M776 606 149 121 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=70050 $D=1
M777 607 149 124 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=74680 $D=1
M778 624 150 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=70050 $D=1
M779 625 150 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=74680 $D=1
M780 151 624 121 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=70050 $D=1
M781 152 625 124 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=74680 $D=1
M782 610 150 151 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=70050 $D=1
M783 611 150 152 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=74680 $D=1
M784 626 153 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=70050 $D=1
M785 627 153 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=74680 $D=1
M786 154 626 151 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=70050 $D=1
M787 155 627 152 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=74680 $D=1
M788 614 153 154 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=70050 $D=1
M789 615 153 155 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=74680 $D=1
M790 628 156 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=70050 $D=1
M791 629 156 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=74680 $D=1
M792 14 628 154 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=70050 $D=1
M793 200 629 155 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=74680 $D=1
M794 618 156 14 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=70050 $D=1
M795 619 156 200 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=74680 $D=1
M796 630 157 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=70050 $D=1
M797 631 157 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=74680 $D=1
M798 632 630 113 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=70050 $D=1
M799 633 631 114 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=74680 $D=1
M800 10 157 632 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=70050 $D=1
M801 11 157 633 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=74680 $D=1
M802 792 539 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=70050 $D=1
M803 793 540 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=74680 $D=1
M804 634 632 792 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=70050 $D=1
M805 635 633 793 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=74680 $D=1
M806 638 539 636 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=70050 $D=1
M807 639 540 637 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=74680 $D=1
M808 636 632 638 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=70050 $D=1
M809 637 633 639 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=74680 $D=1
M810 5 634 636 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=70050 $D=1
M811 6 635 637 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=74680 $D=1
M812 794 640 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=70050 $D=1
M813 795 641 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=74680 $D=1
M814 772 638 794 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=70050 $D=1
M815 773 639 795 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=74680 $D=1
M816 641 772 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=70050 $D=1
M817 158 773 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=74680 $D=1
M818 642 539 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=70050 $D=1
M819 643 540 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=74680 $D=1
M820 5 644 642 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=70050 $D=1
M821 6 645 643 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=74680 $D=1
M822 644 632 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=70050 $D=1
M823 645 633 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=74680 $D=1
M824 796 642 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=70050 $D=1
M825 797 643 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=74680 $D=1
M826 646 640 796 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=70050 $D=1
M827 647 641 797 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=74680 $D=1
M828 649 159 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=70050 $D=1
M829 650 648 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=74680 $D=1
M830 798 646 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=70050 $D=1
M831 799 647 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=74680 $D=1
M832 648 649 798 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=70050 $D=1
M833 160 650 799 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=74680 $D=1
M834 652 651 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=70050 $D=1
M835 653 161 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=74680 $D=1
M836 5 656 654 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=70050 $D=1
M837 6 657 655 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=74680 $D=1
M838 658 116 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=70050 $D=1
M839 659 117 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=74680 $D=1
M840 656 658 651 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=70050 $D=1
M841 657 659 161 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=74680 $D=1
M842 652 116 656 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=70050 $D=1
M843 653 117 657 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=74680 $D=1
M844 660 654 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=70050 $D=1
M845 661 655 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=74680 $D=1
M846 162 660 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=70050 $D=1
M847 651 661 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=74680 $D=1
M848 116 654 162 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=70050 $D=1
M849 117 655 651 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=74680 $D=1
M850 662 162 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=70050 $D=1
M851 663 651 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=74680 $D=1
M852 664 654 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=70050 $D=1
M853 665 655 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=74680 $D=1
M854 201 664 662 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=70050 $D=1
M855 202 665 663 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=74680 $D=1
M856 5 654 201 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=70050 $D=1
M857 6 655 202 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=74680 $D=1
M858 666 163 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=70050 $D=1
M859 667 163 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=74680 $D=1
M860 668 666 201 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=70050 $D=1
M861 669 667 202 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=74680 $D=1
M862 12 163 668 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=70050 $D=1
M863 13 163 669 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=74680 $D=1
M864 670 164 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=70050 $D=1
M865 671 164 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=74680 $D=1
M866 164 670 668 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=70050 $D=1
M867 164 671 669 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=74680 $D=1
M868 5 164 164 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=70050 $D=1
M869 6 164 164 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=74680 $D=1
M870 672 112 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=70050 $D=1
M871 673 112 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=74680 $D=1
M872 5 672 674 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=70050 $D=1
M873 6 673 675 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=74680 $D=1
M874 676 112 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=70050 $D=1
M875 677 112 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=74680 $D=1
M876 678 672 164 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=70050 $D=1
M877 679 673 164 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=74680 $D=1
M878 5 678 774 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=70050 $D=1
M879 6 679 775 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=74680 $D=1
M880 680 774 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=70050 $D=1
M881 681 775 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=74680 $D=1
M882 678 674 680 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=70050 $D=1
M883 679 675 681 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=74680 $D=1
M884 682 112 680 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=70050 $D=1
M885 683 112 681 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=74680 $D=1
M886 5 686 684 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=70050 $D=1
M887 6 687 685 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=74680 $D=1
M888 686 112 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=70050 $D=1
M889 687 112 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=74680 $D=1
M890 776 682 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=70050 $D=1
M891 777 683 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=74680 $D=1
M892 688 684 776 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=70050 $D=1
M893 689 685 777 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=74680 $D=1
M894 5 688 116 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=70050 $D=1
M895 6 689 117 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=74680 $D=1
M896 778 116 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=70050 $D=1
M897 779 117 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=74680 $D=1
M898 688 686 778 5 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=70050 $D=1
M899 689 687 779 6 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=74680 $D=1
M900 176 1 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=71300 $D=0
M901 177 1 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=75930 $D=0
M902 178 1 2 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=71300 $D=0
M903 179 1 3 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=75930 $D=0
M904 5 176 178 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=71300 $D=0
M905 6 177 179 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=75930 $D=0
M906 180 1 4 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=71300 $D=0
M907 181 1 4 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=75930 $D=0
M908 3 176 180 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=71300 $D=0
M909 3 177 181 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=75930 $D=0
M910 182 1 5 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=71300 $D=0
M911 183 1 6 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=75930 $D=0
M912 5 176 182 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=71300 $D=0
M913 3 177 183 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=75930 $D=0
M914 186 7 182 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=71300 $D=0
M915 187 7 183 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=75930 $D=0
M916 184 7 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=71300 $D=0
M917 185 7 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=75930 $D=0
M918 188 7 180 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=71300 $D=0
M919 189 7 181 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=75930 $D=0
M920 178 184 188 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=71300 $D=0
M921 179 185 189 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=75930 $D=0
M922 190 8 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=71300 $D=0
M923 191 8 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=75930 $D=0
M924 192 8 188 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=71300 $D=0
M925 193 8 189 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=75930 $D=0
M926 186 190 192 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=71300 $D=0
M927 187 191 193 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=75930 $D=0
M928 194 9 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=71300 $D=0
M929 195 9 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=75930 $D=0
M930 196 9 5 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=71300 $D=0
M931 197 9 6 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=75930 $D=0
M932 10 194 196 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=71300 $D=0
M933 11 195 197 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=75930 $D=0
M934 198 9 12 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=71300 $D=0
M935 199 9 13 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=75930 $D=0
M936 14 194 198 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=71300 $D=0
M937 200 195 199 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=75930 $D=0
M938 203 9 201 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=71300 $D=0
M939 204 9 202 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=75930 $D=0
M940 192 194 203 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=71300 $D=0
M941 193 195 204 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=75930 $D=0
M942 207 15 203 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=71300 $D=0
M943 208 15 204 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=75930 $D=0
M944 205 15 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=71300 $D=0
M945 206 15 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=75930 $D=0
M946 209 15 198 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=71300 $D=0
M947 210 15 199 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=75930 $D=0
M948 196 205 209 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=71300 $D=0
M949 197 206 210 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=75930 $D=0
M950 211 16 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=71300 $D=0
M951 212 16 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=75930 $D=0
M952 213 16 209 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=71300 $D=0
M953 214 16 210 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=75930 $D=0
M954 207 211 213 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=71300 $D=0
M955 208 212 214 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=75930 $D=0
M956 165 17 215 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=71300 $D=0
M957 166 17 216 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=75930 $D=0
M958 217 18 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=71300 $D=0
M959 218 18 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=75930 $D=0
M960 219 215 213 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=71300 $D=0
M961 220 216 214 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=75930 $D=0
M962 165 219 690 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=71300 $D=0
M963 166 220 691 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=75930 $D=0
M964 221 690 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=71300 $D=0
M965 222 691 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=75930 $D=0
M966 219 17 221 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=71300 $D=0
M967 220 17 222 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=75930 $D=0
M968 221 217 223 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=71300 $D=0
M969 222 218 224 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=75930 $D=0
M970 227 225 221 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=71300 $D=0
M971 228 226 222 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=75930 $D=0
M972 225 19 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=71300 $D=0
M973 226 19 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=75930 $D=0
M974 165 20 229 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=71300 $D=0
M975 166 20 230 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=75930 $D=0
M976 231 21 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=71300 $D=0
M977 232 21 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=75930 $D=0
M978 233 229 213 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=71300 $D=0
M979 234 230 214 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=75930 $D=0
M980 165 233 692 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=71300 $D=0
M981 166 234 693 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=75930 $D=0
M982 235 692 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=71300 $D=0
M983 236 693 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=75930 $D=0
M984 233 20 235 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=71300 $D=0
M985 234 20 236 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=75930 $D=0
M986 235 231 223 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=71300 $D=0
M987 236 232 224 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=75930 $D=0
M988 227 237 235 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=71300 $D=0
M989 228 238 236 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=75930 $D=0
M990 237 22 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=71300 $D=0
M991 238 22 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=75930 $D=0
M992 165 23 239 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=71300 $D=0
M993 166 23 240 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=75930 $D=0
M994 241 24 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=71300 $D=0
M995 242 24 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=75930 $D=0
M996 243 239 213 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=71300 $D=0
M997 244 240 214 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=75930 $D=0
M998 165 243 694 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=71300 $D=0
M999 166 244 695 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=75930 $D=0
M1000 245 694 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=71300 $D=0
M1001 246 695 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=75930 $D=0
M1002 243 23 245 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=71300 $D=0
M1003 244 23 246 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=75930 $D=0
M1004 245 241 223 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=71300 $D=0
M1005 246 242 224 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=75930 $D=0
M1006 227 247 245 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=71300 $D=0
M1007 228 248 246 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=75930 $D=0
M1008 247 25 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=71300 $D=0
M1009 248 25 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=75930 $D=0
M1010 165 26 249 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=71300 $D=0
M1011 166 26 250 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=75930 $D=0
M1012 251 27 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=71300 $D=0
M1013 252 27 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=75930 $D=0
M1014 253 249 213 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=71300 $D=0
M1015 254 250 214 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=75930 $D=0
M1016 165 253 696 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=71300 $D=0
M1017 166 254 697 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=75930 $D=0
M1018 255 696 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=71300 $D=0
M1019 256 697 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=75930 $D=0
M1020 253 26 255 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=71300 $D=0
M1021 254 26 256 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=75930 $D=0
M1022 255 251 223 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=71300 $D=0
M1023 256 252 224 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=75930 $D=0
M1024 227 257 255 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=71300 $D=0
M1025 228 258 256 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=75930 $D=0
M1026 257 28 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=71300 $D=0
M1027 258 28 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=75930 $D=0
M1028 165 29 259 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=71300 $D=0
M1029 166 29 260 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=75930 $D=0
M1030 261 30 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=71300 $D=0
M1031 262 30 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=75930 $D=0
M1032 263 259 213 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=71300 $D=0
M1033 264 260 214 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=75930 $D=0
M1034 165 263 698 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=71300 $D=0
M1035 166 264 699 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=75930 $D=0
M1036 265 698 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=71300 $D=0
M1037 266 699 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=75930 $D=0
M1038 263 29 265 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=71300 $D=0
M1039 264 29 266 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=75930 $D=0
M1040 265 261 223 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=71300 $D=0
M1041 266 262 224 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=75930 $D=0
M1042 227 267 265 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=71300 $D=0
M1043 228 268 266 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=75930 $D=0
M1044 267 31 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=71300 $D=0
M1045 268 31 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=75930 $D=0
M1046 165 32 269 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=71300 $D=0
M1047 166 32 270 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=75930 $D=0
M1048 271 33 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=71300 $D=0
M1049 272 33 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=75930 $D=0
M1050 273 269 213 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=71300 $D=0
M1051 274 270 214 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=75930 $D=0
M1052 165 273 700 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=71300 $D=0
M1053 166 274 701 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=75930 $D=0
M1054 275 700 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=71300 $D=0
M1055 276 701 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=75930 $D=0
M1056 273 32 275 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=71300 $D=0
M1057 274 32 276 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=75930 $D=0
M1058 275 271 223 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=71300 $D=0
M1059 276 272 224 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=75930 $D=0
M1060 227 277 275 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=71300 $D=0
M1061 228 278 276 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=75930 $D=0
M1062 277 34 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=71300 $D=0
M1063 278 34 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=75930 $D=0
M1064 165 35 279 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=71300 $D=0
M1065 166 35 280 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=75930 $D=0
M1066 281 36 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=71300 $D=0
M1067 282 36 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=75930 $D=0
M1068 283 279 213 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=71300 $D=0
M1069 284 280 214 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=75930 $D=0
M1070 165 283 702 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=71300 $D=0
M1071 166 284 703 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=75930 $D=0
M1072 285 702 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=71300 $D=0
M1073 286 703 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=75930 $D=0
M1074 283 35 285 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=71300 $D=0
M1075 284 35 286 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=75930 $D=0
M1076 285 281 223 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=71300 $D=0
M1077 286 282 224 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=75930 $D=0
M1078 227 287 285 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=71300 $D=0
M1079 228 288 286 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=75930 $D=0
M1080 287 37 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=71300 $D=0
M1081 288 37 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=75930 $D=0
M1082 165 38 289 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=71300 $D=0
M1083 166 38 290 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=75930 $D=0
M1084 291 39 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=71300 $D=0
M1085 292 39 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=75930 $D=0
M1086 293 289 213 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=71300 $D=0
M1087 294 290 214 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=75930 $D=0
M1088 165 293 704 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=71300 $D=0
M1089 166 294 705 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=75930 $D=0
M1090 295 704 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=71300 $D=0
M1091 296 705 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=75930 $D=0
M1092 293 38 295 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=71300 $D=0
M1093 294 38 296 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=75930 $D=0
M1094 295 291 223 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=71300 $D=0
M1095 296 292 224 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=75930 $D=0
M1096 227 297 295 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=71300 $D=0
M1097 228 298 296 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=75930 $D=0
M1098 297 40 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=71300 $D=0
M1099 298 40 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=75930 $D=0
M1100 165 41 299 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=71300 $D=0
M1101 166 41 300 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=75930 $D=0
M1102 301 42 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=71300 $D=0
M1103 302 42 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=75930 $D=0
M1104 303 299 213 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=71300 $D=0
M1105 304 300 214 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=75930 $D=0
M1106 165 303 706 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=71300 $D=0
M1107 166 304 707 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=75930 $D=0
M1108 305 706 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=71300 $D=0
M1109 306 707 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=75930 $D=0
M1110 303 41 305 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=71300 $D=0
M1111 304 41 306 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=75930 $D=0
M1112 305 301 223 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=71300 $D=0
M1113 306 302 224 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=75930 $D=0
M1114 227 307 305 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=71300 $D=0
M1115 228 308 306 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=75930 $D=0
M1116 307 43 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=71300 $D=0
M1117 308 43 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=75930 $D=0
M1118 165 44 309 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=71300 $D=0
M1119 166 44 310 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=75930 $D=0
M1120 311 45 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=71300 $D=0
M1121 312 45 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=75930 $D=0
M1122 313 309 213 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=71300 $D=0
M1123 314 310 214 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=75930 $D=0
M1124 165 313 708 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=71300 $D=0
M1125 166 314 709 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=75930 $D=0
M1126 315 708 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=71300 $D=0
M1127 316 709 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=75930 $D=0
M1128 313 44 315 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=71300 $D=0
M1129 314 44 316 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=75930 $D=0
M1130 315 311 223 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=71300 $D=0
M1131 316 312 224 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=75930 $D=0
M1132 227 317 315 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=71300 $D=0
M1133 228 318 316 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=75930 $D=0
M1134 317 46 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=71300 $D=0
M1135 318 46 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=75930 $D=0
M1136 165 47 319 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=71300 $D=0
M1137 166 47 320 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=75930 $D=0
M1138 321 48 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=71300 $D=0
M1139 322 48 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=75930 $D=0
M1140 323 319 213 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=71300 $D=0
M1141 324 320 214 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=75930 $D=0
M1142 165 323 710 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=71300 $D=0
M1143 166 324 711 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=75930 $D=0
M1144 325 710 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=71300 $D=0
M1145 326 711 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=75930 $D=0
M1146 323 47 325 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=71300 $D=0
M1147 324 47 326 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=75930 $D=0
M1148 325 321 223 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=71300 $D=0
M1149 326 322 224 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=75930 $D=0
M1150 227 327 325 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=71300 $D=0
M1151 228 328 326 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=75930 $D=0
M1152 327 49 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=71300 $D=0
M1153 328 49 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=75930 $D=0
M1154 165 50 329 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=71300 $D=0
M1155 166 50 330 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=75930 $D=0
M1156 331 51 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=71300 $D=0
M1157 332 51 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=75930 $D=0
M1158 333 329 213 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=71300 $D=0
M1159 334 330 214 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=75930 $D=0
M1160 165 333 712 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=71300 $D=0
M1161 166 334 713 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=75930 $D=0
M1162 335 712 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=71300 $D=0
M1163 336 713 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=75930 $D=0
M1164 333 50 335 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=71300 $D=0
M1165 334 50 336 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=75930 $D=0
M1166 335 331 223 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=71300 $D=0
M1167 336 332 224 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=75930 $D=0
M1168 227 337 335 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=71300 $D=0
M1169 228 338 336 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=75930 $D=0
M1170 337 52 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=71300 $D=0
M1171 338 52 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=75930 $D=0
M1172 165 53 339 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=71300 $D=0
M1173 166 53 340 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=75930 $D=0
M1174 341 54 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=71300 $D=0
M1175 342 54 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=75930 $D=0
M1176 343 339 213 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=71300 $D=0
M1177 344 340 214 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=75930 $D=0
M1178 165 343 714 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=71300 $D=0
M1179 166 344 715 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=75930 $D=0
M1180 345 714 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=71300 $D=0
M1181 346 715 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=75930 $D=0
M1182 343 53 345 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=71300 $D=0
M1183 344 53 346 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=75930 $D=0
M1184 345 341 223 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=71300 $D=0
M1185 346 342 224 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=75930 $D=0
M1186 227 347 345 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=71300 $D=0
M1187 228 348 346 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=75930 $D=0
M1188 347 55 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=71300 $D=0
M1189 348 55 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=75930 $D=0
M1190 165 56 349 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=71300 $D=0
M1191 166 56 350 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=75930 $D=0
M1192 351 57 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=71300 $D=0
M1193 352 57 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=75930 $D=0
M1194 353 349 213 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=71300 $D=0
M1195 354 350 214 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=75930 $D=0
M1196 165 353 716 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=71300 $D=0
M1197 166 354 717 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=75930 $D=0
M1198 355 716 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=71300 $D=0
M1199 356 717 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=75930 $D=0
M1200 353 56 355 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=71300 $D=0
M1201 354 56 356 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=75930 $D=0
M1202 355 351 223 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=71300 $D=0
M1203 356 352 224 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=75930 $D=0
M1204 227 357 355 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=71300 $D=0
M1205 228 358 356 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=75930 $D=0
M1206 357 58 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=71300 $D=0
M1207 358 58 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=75930 $D=0
M1208 165 59 359 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=71300 $D=0
M1209 166 59 360 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=75930 $D=0
M1210 361 60 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=71300 $D=0
M1211 362 60 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=75930 $D=0
M1212 363 359 213 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=71300 $D=0
M1213 364 360 214 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=75930 $D=0
M1214 165 363 718 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=71300 $D=0
M1215 166 364 719 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=75930 $D=0
M1216 365 718 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=71300 $D=0
M1217 366 719 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=75930 $D=0
M1218 363 59 365 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=71300 $D=0
M1219 364 59 366 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=75930 $D=0
M1220 365 361 223 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=71300 $D=0
M1221 366 362 224 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=75930 $D=0
M1222 227 367 365 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=71300 $D=0
M1223 228 368 366 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=75930 $D=0
M1224 367 61 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=71300 $D=0
M1225 368 61 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=75930 $D=0
M1226 165 62 369 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=71300 $D=0
M1227 166 62 370 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=75930 $D=0
M1228 371 63 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=71300 $D=0
M1229 372 63 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=75930 $D=0
M1230 373 369 213 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=71300 $D=0
M1231 374 370 214 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=75930 $D=0
M1232 165 373 720 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=71300 $D=0
M1233 166 374 721 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=75930 $D=0
M1234 375 720 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=71300 $D=0
M1235 376 721 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=75930 $D=0
M1236 373 62 375 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=71300 $D=0
M1237 374 62 376 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=75930 $D=0
M1238 375 371 223 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=71300 $D=0
M1239 376 372 224 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=75930 $D=0
M1240 227 377 375 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=71300 $D=0
M1241 228 378 376 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=75930 $D=0
M1242 377 64 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=71300 $D=0
M1243 378 64 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=75930 $D=0
M1244 165 65 379 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=71300 $D=0
M1245 166 65 380 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=75930 $D=0
M1246 381 66 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=71300 $D=0
M1247 382 66 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=75930 $D=0
M1248 383 379 213 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=71300 $D=0
M1249 384 380 214 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=75930 $D=0
M1250 165 383 722 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=71300 $D=0
M1251 166 384 723 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=75930 $D=0
M1252 385 722 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=71300 $D=0
M1253 386 723 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=75930 $D=0
M1254 383 65 385 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=71300 $D=0
M1255 384 65 386 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=75930 $D=0
M1256 385 381 223 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=71300 $D=0
M1257 386 382 224 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=75930 $D=0
M1258 227 387 385 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=71300 $D=0
M1259 228 388 386 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=75930 $D=0
M1260 387 67 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=71300 $D=0
M1261 388 67 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=75930 $D=0
M1262 165 68 389 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=71300 $D=0
M1263 166 68 390 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=75930 $D=0
M1264 391 69 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=71300 $D=0
M1265 392 69 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=75930 $D=0
M1266 393 389 213 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=71300 $D=0
M1267 394 390 214 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=75930 $D=0
M1268 165 393 724 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=71300 $D=0
M1269 166 394 725 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=75930 $D=0
M1270 395 724 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=71300 $D=0
M1271 396 725 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=75930 $D=0
M1272 393 68 395 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=71300 $D=0
M1273 394 68 396 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=75930 $D=0
M1274 395 391 223 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=71300 $D=0
M1275 396 392 224 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=75930 $D=0
M1276 227 397 395 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=71300 $D=0
M1277 228 398 396 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=75930 $D=0
M1278 397 70 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=71300 $D=0
M1279 398 70 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=75930 $D=0
M1280 165 71 399 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=71300 $D=0
M1281 166 71 400 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=75930 $D=0
M1282 401 72 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=71300 $D=0
M1283 402 72 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=75930 $D=0
M1284 403 399 213 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=71300 $D=0
M1285 404 400 214 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=75930 $D=0
M1286 165 403 726 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=71300 $D=0
M1287 166 404 727 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=75930 $D=0
M1288 405 726 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=71300 $D=0
M1289 406 727 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=75930 $D=0
M1290 403 71 405 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=71300 $D=0
M1291 404 71 406 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=75930 $D=0
M1292 405 401 223 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=71300 $D=0
M1293 406 402 224 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=75930 $D=0
M1294 227 407 405 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=71300 $D=0
M1295 228 408 406 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=75930 $D=0
M1296 407 73 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=71300 $D=0
M1297 408 73 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=75930 $D=0
M1298 165 74 409 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=71300 $D=0
M1299 166 74 410 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=75930 $D=0
M1300 411 75 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=71300 $D=0
M1301 412 75 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=75930 $D=0
M1302 413 409 213 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=71300 $D=0
M1303 414 410 214 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=75930 $D=0
M1304 165 413 728 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=71300 $D=0
M1305 166 414 729 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=75930 $D=0
M1306 415 728 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=71300 $D=0
M1307 416 729 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=75930 $D=0
M1308 413 74 415 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=71300 $D=0
M1309 414 74 416 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=75930 $D=0
M1310 415 411 223 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=71300 $D=0
M1311 416 412 224 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=75930 $D=0
M1312 227 417 415 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=71300 $D=0
M1313 228 418 416 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=75930 $D=0
M1314 417 76 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=71300 $D=0
M1315 418 76 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=75930 $D=0
M1316 165 77 419 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=71300 $D=0
M1317 166 77 420 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=75930 $D=0
M1318 421 78 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=71300 $D=0
M1319 422 78 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=75930 $D=0
M1320 423 419 213 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=71300 $D=0
M1321 424 420 214 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=75930 $D=0
M1322 165 423 730 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=71300 $D=0
M1323 166 424 731 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=75930 $D=0
M1324 425 730 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=71300 $D=0
M1325 426 731 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=75930 $D=0
M1326 423 77 425 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=71300 $D=0
M1327 424 77 426 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=75930 $D=0
M1328 425 421 223 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=71300 $D=0
M1329 426 422 224 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=75930 $D=0
M1330 227 427 425 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=71300 $D=0
M1331 228 428 426 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=75930 $D=0
M1332 427 79 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=71300 $D=0
M1333 428 79 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=75930 $D=0
M1334 165 80 429 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=71300 $D=0
M1335 166 80 430 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=75930 $D=0
M1336 431 81 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=71300 $D=0
M1337 432 81 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=75930 $D=0
M1338 433 429 213 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=71300 $D=0
M1339 434 430 214 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=75930 $D=0
M1340 165 433 732 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=71300 $D=0
M1341 166 434 733 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=75930 $D=0
M1342 435 732 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=71300 $D=0
M1343 436 733 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=75930 $D=0
M1344 433 80 435 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=71300 $D=0
M1345 434 80 436 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=75930 $D=0
M1346 435 431 223 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=71300 $D=0
M1347 436 432 224 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=75930 $D=0
M1348 227 437 435 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=71300 $D=0
M1349 228 438 436 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=75930 $D=0
M1350 437 82 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=71300 $D=0
M1351 438 82 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=75930 $D=0
M1352 165 83 439 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=71300 $D=0
M1353 166 83 440 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=75930 $D=0
M1354 441 84 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=71300 $D=0
M1355 442 84 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=75930 $D=0
M1356 443 439 213 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=71300 $D=0
M1357 444 440 214 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=75930 $D=0
M1358 165 443 734 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=71300 $D=0
M1359 166 444 735 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=75930 $D=0
M1360 445 734 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=71300 $D=0
M1361 446 735 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=75930 $D=0
M1362 443 83 445 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=71300 $D=0
M1363 444 83 446 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=75930 $D=0
M1364 445 441 223 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=71300 $D=0
M1365 446 442 224 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=75930 $D=0
M1366 227 447 445 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=71300 $D=0
M1367 228 448 446 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=75930 $D=0
M1368 447 85 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=71300 $D=0
M1369 448 85 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=75930 $D=0
M1370 165 86 449 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=71300 $D=0
M1371 166 86 450 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=75930 $D=0
M1372 451 87 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=71300 $D=0
M1373 452 87 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=75930 $D=0
M1374 453 449 213 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=71300 $D=0
M1375 454 450 214 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=75930 $D=0
M1376 165 453 736 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=71300 $D=0
M1377 166 454 737 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=75930 $D=0
M1378 455 736 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=71300 $D=0
M1379 456 737 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=75930 $D=0
M1380 453 86 455 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=71300 $D=0
M1381 454 86 456 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=75930 $D=0
M1382 455 451 223 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=71300 $D=0
M1383 456 452 224 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=75930 $D=0
M1384 227 457 455 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=71300 $D=0
M1385 228 458 456 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=75930 $D=0
M1386 457 88 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=71300 $D=0
M1387 458 88 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=75930 $D=0
M1388 165 89 459 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=71300 $D=0
M1389 166 89 460 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=75930 $D=0
M1390 461 90 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=71300 $D=0
M1391 462 90 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=75930 $D=0
M1392 463 459 213 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=71300 $D=0
M1393 464 460 214 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=75930 $D=0
M1394 165 463 738 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=71300 $D=0
M1395 166 464 739 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=75930 $D=0
M1396 465 738 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=71300 $D=0
M1397 466 739 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=75930 $D=0
M1398 463 89 465 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=71300 $D=0
M1399 464 89 466 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=75930 $D=0
M1400 465 461 223 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=71300 $D=0
M1401 466 462 224 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=75930 $D=0
M1402 227 467 465 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=71300 $D=0
M1403 228 468 466 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=75930 $D=0
M1404 467 91 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=71300 $D=0
M1405 468 91 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=75930 $D=0
M1406 165 92 469 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=71300 $D=0
M1407 166 92 470 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=75930 $D=0
M1408 471 93 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=71300 $D=0
M1409 472 93 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=75930 $D=0
M1410 473 469 213 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=71300 $D=0
M1411 474 470 214 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=75930 $D=0
M1412 165 473 740 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=71300 $D=0
M1413 166 474 741 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=75930 $D=0
M1414 475 740 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=71300 $D=0
M1415 476 741 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=75930 $D=0
M1416 473 92 475 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=71300 $D=0
M1417 474 92 476 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=75930 $D=0
M1418 475 471 223 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=71300 $D=0
M1419 476 472 224 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=75930 $D=0
M1420 227 477 475 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=71300 $D=0
M1421 228 478 476 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=75930 $D=0
M1422 477 94 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=71300 $D=0
M1423 478 94 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=75930 $D=0
M1424 165 95 479 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=71300 $D=0
M1425 166 95 480 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=75930 $D=0
M1426 481 96 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=71300 $D=0
M1427 482 96 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=75930 $D=0
M1428 483 479 213 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=71300 $D=0
M1429 484 480 214 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=75930 $D=0
M1430 165 483 742 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=71300 $D=0
M1431 166 484 743 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=75930 $D=0
M1432 485 742 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=71300 $D=0
M1433 486 743 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=75930 $D=0
M1434 483 95 485 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=71300 $D=0
M1435 484 95 486 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=75930 $D=0
M1436 485 481 223 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=71300 $D=0
M1437 486 482 224 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=75930 $D=0
M1438 227 487 485 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=71300 $D=0
M1439 228 488 486 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=75930 $D=0
M1440 487 97 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=71300 $D=0
M1441 488 97 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=75930 $D=0
M1442 165 98 489 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=71300 $D=0
M1443 166 98 490 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=75930 $D=0
M1444 491 99 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=71300 $D=0
M1445 492 99 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=75930 $D=0
M1446 493 489 213 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=71300 $D=0
M1447 494 490 214 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=75930 $D=0
M1448 165 493 744 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=71300 $D=0
M1449 166 494 745 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=75930 $D=0
M1450 495 744 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=71300 $D=0
M1451 496 745 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=75930 $D=0
M1452 493 98 495 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=71300 $D=0
M1453 494 98 496 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=75930 $D=0
M1454 495 491 223 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=71300 $D=0
M1455 496 492 224 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=75930 $D=0
M1456 227 497 495 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=71300 $D=0
M1457 228 498 496 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=75930 $D=0
M1458 497 100 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=71300 $D=0
M1459 498 100 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=75930 $D=0
M1460 165 101 499 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=71300 $D=0
M1461 166 101 500 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=75930 $D=0
M1462 501 102 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=71300 $D=0
M1463 502 102 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=75930 $D=0
M1464 503 499 213 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=71300 $D=0
M1465 504 500 214 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=75930 $D=0
M1466 165 503 746 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=71300 $D=0
M1467 166 504 747 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=75930 $D=0
M1468 505 746 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=71300 $D=0
M1469 506 747 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=75930 $D=0
M1470 503 101 505 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=71300 $D=0
M1471 504 101 506 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=75930 $D=0
M1472 505 501 223 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=71300 $D=0
M1473 506 502 224 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=75930 $D=0
M1474 227 507 505 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=71300 $D=0
M1475 228 508 506 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=75930 $D=0
M1476 507 103 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=71300 $D=0
M1477 508 103 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=75930 $D=0
M1478 165 104 509 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=71300 $D=0
M1479 166 104 510 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=75930 $D=0
M1480 511 105 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=71300 $D=0
M1481 512 105 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=75930 $D=0
M1482 513 509 213 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=71300 $D=0
M1483 514 510 214 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=75930 $D=0
M1484 165 513 748 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=71300 $D=0
M1485 166 514 749 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=75930 $D=0
M1486 515 748 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=71300 $D=0
M1487 516 749 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=75930 $D=0
M1488 513 104 515 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=71300 $D=0
M1489 514 104 516 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=75930 $D=0
M1490 515 511 223 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=71300 $D=0
M1491 516 512 224 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=75930 $D=0
M1492 227 517 515 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=71300 $D=0
M1493 228 518 516 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=75930 $D=0
M1494 517 106 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=71300 $D=0
M1495 518 106 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=75930 $D=0
M1496 165 107 519 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=71300 $D=0
M1497 166 107 520 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=75930 $D=0
M1498 521 108 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=71300 $D=0
M1499 522 108 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=75930 $D=0
M1500 523 519 213 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=71300 $D=0
M1501 524 520 214 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=75930 $D=0
M1502 165 523 750 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=71300 $D=0
M1503 166 524 751 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=75930 $D=0
M1504 525 750 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=71300 $D=0
M1505 526 751 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=75930 $D=0
M1506 523 107 525 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=71300 $D=0
M1507 524 107 526 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=75930 $D=0
M1508 525 521 223 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=71300 $D=0
M1509 526 522 224 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=75930 $D=0
M1510 227 527 525 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=71300 $D=0
M1511 228 528 526 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=75930 $D=0
M1512 527 109 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=71300 $D=0
M1513 528 109 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=75930 $D=0
M1514 165 110 529 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=71300 $D=0
M1515 166 110 530 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=75930 $D=0
M1516 531 111 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=71300 $D=0
M1517 532 111 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=75930 $D=0
M1518 5 531 223 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=71300 $D=0
M1519 6 532 224 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=75930 $D=0
M1520 227 529 5 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=71300 $D=0
M1521 228 530 6 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=75930 $D=0
M1522 165 535 533 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=71300 $D=0
M1523 166 536 534 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=75930 $D=0
M1524 535 112 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=71300 $D=0
M1525 536 112 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=75930 $D=0
M1526 752 223 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=71300 $D=0
M1527 753 224 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=75930 $D=0
M1528 537 535 752 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=71300 $D=0
M1529 538 536 753 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=75930 $D=0
M1530 165 537 539 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=71300 $D=0
M1531 166 538 540 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=75930 $D=0
M1532 754 539 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=71300 $D=0
M1533 755 540 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=75930 $D=0
M1534 537 533 754 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=71300 $D=0
M1535 538 534 755 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=75930 $D=0
M1536 165 543 541 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=71300 $D=0
M1537 166 544 542 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=75930 $D=0
M1538 543 112 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=71300 $D=0
M1539 544 112 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=75930 $D=0
M1540 756 227 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=71300 $D=0
M1541 757 228 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=75930 $D=0
M1542 545 543 756 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=71300 $D=0
M1543 546 544 757 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=75930 $D=0
M1544 165 545 113 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=71300 $D=0
M1545 166 546 114 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=75930 $D=0
M1546 758 113 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=71300 $D=0
M1547 759 114 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=75930 $D=0
M1548 545 541 758 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=71300 $D=0
M1549 546 542 759 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=75930 $D=0
M1550 547 115 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=71300 $D=0
M1551 548 115 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=75930 $D=0
M1552 549 115 539 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=71300 $D=0
M1553 550 115 540 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=75930 $D=0
M1554 116 547 549 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=71300 $D=0
M1555 117 548 550 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=75930 $D=0
M1556 551 118 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=71300 $D=0
M1557 552 118 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=75930 $D=0
M1558 553 118 113 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=71300 $D=0
M1559 554 118 114 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=75930 $D=0
M1560 760 551 553 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=71300 $D=0
M1561 761 552 554 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=75930 $D=0
M1562 165 113 760 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=71300 $D=0
M1563 166 114 761 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=75930 $D=0
M1564 555 119 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=71300 $D=0
M1565 556 119 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=75930 $D=0
M1566 557 119 553 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=71300 $D=0
M1567 558 119 554 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=75930 $D=0
M1568 10 555 557 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=71300 $D=0
M1569 11 556 558 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=75930 $D=0
M1570 560 559 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=71300 $D=0
M1571 561 120 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=75930 $D=0
M1572 165 564 562 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=71300 $D=0
M1573 166 565 563 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=75930 $D=0
M1574 566 549 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=71300 $D=0
M1575 567 550 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=75930 $D=0
M1576 564 549 559 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=71300 $D=0
M1577 565 550 120 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=75930 $D=0
M1578 560 566 564 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=71300 $D=0
M1579 561 567 565 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=75930 $D=0
M1580 568 562 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=71300 $D=0
M1581 569 563 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=75930 $D=0
M1582 570 562 557 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=71300 $D=0
M1583 559 563 558 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=75930 $D=0
M1584 549 568 570 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=71300 $D=0
M1585 550 569 559 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=75930 $D=0
M1586 571 570 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=71300 $D=0
M1587 572 559 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=75930 $D=0
M1588 573 562 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=71300 $D=0
M1589 574 563 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=75930 $D=0
M1590 575 562 571 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=71300 $D=0
M1591 576 563 572 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=75930 $D=0
M1592 557 573 575 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=71300 $D=0
M1593 558 574 576 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=75930 $D=0
M1594 780 549 165 165 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=70940 $D=0
M1595 781 550 166 166 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=75570 $D=0
M1596 577 557 780 165 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=70940 $D=0
M1597 578 558 781 166 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=75570 $D=0
M1598 579 575 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=71300 $D=0
M1599 580 576 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=75930 $D=0
M1600 581 549 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=71300 $D=0
M1601 582 550 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=75930 $D=0
M1602 165 557 581 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=71300 $D=0
M1603 166 558 582 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=75930 $D=0
M1604 583 549 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=71300 $D=0
M1605 584 550 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=75930 $D=0
M1606 165 557 583 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=71300 $D=0
M1607 166 558 584 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=75930 $D=0
M1608 782 549 165 165 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=71120 $D=0
M1609 783 550 166 166 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=75750 $D=0
M1610 587 557 782 165 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=71120 $D=0
M1611 588 558 783 166 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=75750 $D=0
M1612 165 583 587 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=71300 $D=0
M1613 166 584 588 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=75930 $D=0
M1614 589 125 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=71300 $D=0
M1615 590 125 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=75930 $D=0
M1616 591 125 577 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=71300 $D=0
M1617 592 125 578 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=75930 $D=0
M1618 581 589 591 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=71300 $D=0
M1619 582 590 592 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=75930 $D=0
M1620 593 125 579 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=71300 $D=0
M1621 594 125 580 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=75930 $D=0
M1622 587 589 593 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=71300 $D=0
M1623 588 590 594 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=75930 $D=0
M1624 595 126 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=71300 $D=0
M1625 596 126 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=75930 $D=0
M1626 597 126 593 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=71300 $D=0
M1627 598 126 594 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=75930 $D=0
M1628 591 595 597 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=71300 $D=0
M1629 592 596 598 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=75930 $D=0
M1630 12 597 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=71300 $D=0
M1631 13 598 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=75930 $D=0
M1632 599 127 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=71300 $D=0
M1633 600 127 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=75930 $D=0
M1634 601 127 128 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=71300 $D=0
M1635 602 127 129 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=75930 $D=0
M1636 130 599 601 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=71300 $D=0
M1637 131 600 602 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=75930 $D=0
M1638 603 127 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=71300 $D=0
M1639 604 127 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=75930 $D=0
M1640 606 127 132 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=71300 $D=0
M1641 607 127 133 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=75930 $D=0
M1642 134 603 606 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=71300 $D=0
M1643 135 604 607 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=75930 $D=0
M1644 608 127 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=71300 $D=0
M1645 609 127 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=75930 $D=0
M1646 610 127 122 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=71300 $D=0
M1647 611 127 136 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=75930 $D=0
M1648 137 608 610 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=71300 $D=0
M1649 138 609 611 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=75930 $D=0
M1650 612 127 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=71300 $D=0
M1651 613 127 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=75930 $D=0
M1652 614 127 139 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=71300 $D=0
M1653 615 127 140 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=75930 $D=0
M1654 141 612 614 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=71300 $D=0
M1655 142 613 615 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=75930 $D=0
M1656 616 127 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=71300 $D=0
M1657 617 127 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=75930 $D=0
M1658 618 127 143 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=71300 $D=0
M1659 619 127 6 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=75930 $D=0
M1660 144 616 618 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=71300 $D=0
M1661 145 617 619 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=75930 $D=0
M1662 165 549 770 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=71300 $D=0
M1663 166 550 771 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=75930 $D=0
M1664 131 770 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=71300 $D=0
M1665 128 771 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=75930 $D=0
M1666 620 146 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=71300 $D=0
M1667 621 146 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=75930 $D=0
M1668 147 146 131 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=71300 $D=0
M1669 148 146 128 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=75930 $D=0
M1670 601 620 147 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=71300 $D=0
M1671 602 621 148 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=75930 $D=0
M1672 622 149 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=71300 $D=0
M1673 623 149 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=75930 $D=0
M1674 121 149 147 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=71300 $D=0
M1675 124 149 148 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=75930 $D=0
M1676 606 622 121 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=71300 $D=0
M1677 607 623 124 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=75930 $D=0
M1678 624 150 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=71300 $D=0
M1679 625 150 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=75930 $D=0
M1680 151 150 121 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=71300 $D=0
M1681 152 150 124 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=75930 $D=0
M1682 610 624 151 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=71300 $D=0
M1683 611 625 152 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=75930 $D=0
M1684 626 153 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=71300 $D=0
M1685 627 153 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=75930 $D=0
M1686 154 153 151 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=71300 $D=0
M1687 155 153 152 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=75930 $D=0
M1688 614 626 154 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=71300 $D=0
M1689 615 627 155 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=75930 $D=0
M1690 628 156 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=71300 $D=0
M1691 629 156 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=75930 $D=0
M1692 14 156 154 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=71300 $D=0
M1693 200 156 155 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=75930 $D=0
M1694 618 628 14 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=71300 $D=0
M1695 619 629 200 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=75930 $D=0
M1696 630 157 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=71300 $D=0
M1697 631 157 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=75930 $D=0
M1698 632 157 113 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=71300 $D=0
M1699 633 157 114 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=75930 $D=0
M1700 10 630 632 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=71300 $D=0
M1701 11 631 633 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=75930 $D=0
M1702 634 539 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=71300 $D=0
M1703 635 540 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=75930 $D=0
M1704 165 632 634 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=71300 $D=0
M1705 166 633 635 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=75930 $D=0
M1706 784 539 165 165 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=71120 $D=0
M1707 785 540 166 166 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=75750 $D=0
M1708 638 632 784 165 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=71120 $D=0
M1709 639 633 785 166 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=75750 $D=0
M1710 165 634 638 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=71300 $D=0
M1711 166 635 639 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=75930 $D=0
M1712 772 640 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=71300 $D=0
M1713 773 641 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=75930 $D=0
M1714 165 638 772 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=71300 $D=0
M1715 166 639 773 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=75930 $D=0
M1716 641 772 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=71300 $D=0
M1717 158 773 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=75930 $D=0
M1718 786 539 165 165 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=70940 $D=0
M1719 787 540 166 166 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=75570 $D=0
M1720 642 644 786 165 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=70940 $D=0
M1721 643 645 787 166 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=75570 $D=0
M1722 644 632 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=71300 $D=0
M1723 645 633 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=75930 $D=0
M1724 646 642 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=71300 $D=0
M1725 647 643 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=75930 $D=0
M1726 165 640 646 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=71300 $D=0
M1727 166 641 647 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=75930 $D=0
M1728 649 159 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=71300 $D=0
M1729 650 648 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=75930 $D=0
M1730 648 646 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=71300 $D=0
M1731 160 647 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=75930 $D=0
M1732 165 649 648 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=71300 $D=0
M1733 166 650 160 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=75930 $D=0
M1734 652 651 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=71300 $D=0
M1735 653 161 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=75930 $D=0
M1736 165 656 654 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=71300 $D=0
M1737 166 657 655 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=75930 $D=0
M1738 658 116 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=71300 $D=0
M1739 659 117 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=75930 $D=0
M1740 656 116 651 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=71300 $D=0
M1741 657 117 161 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=75930 $D=0
M1742 652 658 656 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=71300 $D=0
M1743 653 659 657 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=75930 $D=0
M1744 660 654 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=71300 $D=0
M1745 661 655 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=75930 $D=0
M1746 162 654 5 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=71300 $D=0
M1747 651 655 6 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=75930 $D=0
M1748 116 660 162 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=71300 $D=0
M1749 117 661 651 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=75930 $D=0
M1750 662 162 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=71300 $D=0
M1751 663 651 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=75930 $D=0
M1752 664 654 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=71300 $D=0
M1753 665 655 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=75930 $D=0
M1754 201 654 662 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=71300 $D=0
M1755 202 655 663 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=75930 $D=0
M1756 5 664 201 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=71300 $D=0
M1757 6 665 202 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=75930 $D=0
M1758 666 163 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=71300 $D=0
M1759 667 163 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=75930 $D=0
M1760 668 163 201 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=71300 $D=0
M1761 669 163 202 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=75930 $D=0
M1762 12 666 668 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=71300 $D=0
M1763 13 667 669 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=75930 $D=0
M1764 670 164 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=71300 $D=0
M1765 671 164 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=75930 $D=0
M1766 164 164 668 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=71300 $D=0
M1767 164 164 669 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=75930 $D=0
M1768 5 670 164 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=71300 $D=0
M1769 6 671 164 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=75930 $D=0
M1770 672 112 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=71300 $D=0
M1771 673 112 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=75930 $D=0
M1772 165 672 674 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=71300 $D=0
M1773 166 673 675 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=75930 $D=0
M1774 676 112 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=71300 $D=0
M1775 677 112 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=75930 $D=0
M1776 678 674 164 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=71300 $D=0
M1777 679 675 164 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=75930 $D=0
M1778 165 678 774 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=71300 $D=0
M1779 166 679 775 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=75930 $D=0
M1780 680 774 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=71300 $D=0
M1781 681 775 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=75930 $D=0
M1782 678 672 680 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=71300 $D=0
M1783 679 673 681 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=75930 $D=0
M1784 682 676 680 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=71300 $D=0
M1785 683 677 681 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=75930 $D=0
M1786 165 686 684 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=71300 $D=0
M1787 166 687 685 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=75930 $D=0
M1788 686 112 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=71300 $D=0
M1789 687 112 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=75930 $D=0
M1790 776 682 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=71300 $D=0
M1791 777 683 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=75930 $D=0
M1792 688 686 776 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=71300 $D=0
M1793 689 687 777 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=75930 $D=0
M1794 165 688 116 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=71300 $D=0
M1795 166 689 117 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=75930 $D=0
M1796 778 116 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=71300 $D=0
M1797 779 117 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=75930 $D=0
M1798 688 684 778 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=71300 $D=0
M1799 689 685 779 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=75930 $D=0
.ENDS
***************************************
.SUBCKT ICV_32
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_33
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_34
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_35
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_36 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180
+ 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200
+ 201 202 203 204 205
** N=1449 EP=205 IP=2964 FDC=3600
M0 208 1 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=51530 $D=1
M1 209 1 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=56160 $D=1
M2 210 1 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=60790 $D=1
M3 211 1 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=65420 $D=1
M4 212 208 2 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=51530 $D=1
M5 213 209 3 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=56160 $D=1
M6 214 210 4 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=60790 $D=1
M7 215 211 5 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=65420 $D=1
M8 8 1 212 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=51530 $D=1
M9 9 1 213 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=56160 $D=1
M10 10 1 214 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=60790 $D=1
M11 11 1 215 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=65420 $D=1
M12 216 208 6 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=51530 $D=1
M13 217 209 6 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=56160 $D=1
M14 218 210 6 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=60790 $D=1
M15 219 211 6 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=65420 $D=1
M16 7 1 216 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=51530 $D=1
M17 7 1 217 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=56160 $D=1
M18 7 1 218 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=60790 $D=1
M19 7 1 219 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=65420 $D=1
M20 220 208 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=51530 $D=1
M21 221 209 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=56160 $D=1
M22 222 210 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=60790 $D=1
M23 223 211 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=65420 $D=1
M24 8 1 220 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=51530 $D=1
M25 9 1 221 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=56160 $D=1
M26 10 1 222 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=60790 $D=1
M27 11 1 223 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=65420 $D=1
M28 228 224 220 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=51530 $D=1
M29 229 225 221 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=56160 $D=1
M30 230 226 222 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=60790 $D=1
M31 231 227 223 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=65420 $D=1
M32 224 12 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=51530 $D=1
M33 225 12 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=56160 $D=1
M34 226 12 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=60790 $D=1
M35 227 12 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=65420 $D=1
M36 232 224 216 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=51530 $D=1
M37 233 225 217 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=56160 $D=1
M38 234 226 218 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=60790 $D=1
M39 235 227 219 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=65420 $D=1
M40 212 12 232 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=51530 $D=1
M41 213 12 233 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=56160 $D=1
M42 214 12 234 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=60790 $D=1
M43 215 12 235 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=65420 $D=1
M44 236 13 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=51530 $D=1
M45 237 13 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=56160 $D=1
M46 238 13 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=60790 $D=1
M47 239 13 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=65420 $D=1
M48 240 236 232 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=51530 $D=1
M49 241 237 233 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=56160 $D=1
M50 242 238 234 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=60790 $D=1
M51 243 239 235 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=65420 $D=1
M52 228 13 240 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=51530 $D=1
M53 229 13 241 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=56160 $D=1
M54 230 13 242 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=60790 $D=1
M55 231 13 243 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=65420 $D=1
M56 244 14 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=51530 $D=1
M57 245 14 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=56160 $D=1
M58 246 14 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=60790 $D=1
M59 247 14 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=65420 $D=1
M60 248 244 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=51530 $D=1
M61 249 245 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=56160 $D=1
M62 250 246 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=60790 $D=1
M63 251 247 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=65420 $D=1
M64 15 14 248 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=51530 $D=1
M65 16 14 249 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=56160 $D=1
M66 17 14 250 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=60790 $D=1
M67 18 14 251 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=65420 $D=1
M68 252 244 19 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=51530 $D=1
M69 253 245 20 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=56160 $D=1
M70 254 246 21 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=60790 $D=1
M71 255 247 22 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=65420 $D=1
M72 23 14 252 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=51530 $D=1
M73 24 14 253 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=56160 $D=1
M74 25 14 254 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=60790 $D=1
M75 26 14 255 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=65420 $D=1
M76 260 244 256 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=51530 $D=1
M77 261 245 257 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=56160 $D=1
M78 262 246 258 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=60790 $D=1
M79 263 247 259 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=65420 $D=1
M80 240 14 260 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=51530 $D=1
M81 241 14 261 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=56160 $D=1
M82 242 14 262 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=60790 $D=1
M83 243 14 263 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=65420 $D=1
M84 268 264 260 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=51530 $D=1
M85 269 265 261 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=56160 $D=1
M86 270 266 262 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=60790 $D=1
M87 271 267 263 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=65420 $D=1
M88 264 27 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=51530 $D=1
M89 265 27 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=56160 $D=1
M90 266 27 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=60790 $D=1
M91 267 27 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=65420 $D=1
M92 272 264 252 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=51530 $D=1
M93 273 265 253 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=56160 $D=1
M94 274 266 254 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=60790 $D=1
M95 275 267 255 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=65420 $D=1
M96 248 27 272 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=51530 $D=1
M97 249 27 273 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=56160 $D=1
M98 250 27 274 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=60790 $D=1
M99 251 27 275 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=65420 $D=1
M100 276 28 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=51530 $D=1
M101 277 28 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=56160 $D=1
M102 278 28 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=60790 $D=1
M103 279 28 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=65420 $D=1
M104 280 276 272 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=51530 $D=1
M105 281 277 273 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=56160 $D=1
M106 282 278 274 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=60790 $D=1
M107 283 279 275 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=65420 $D=1
M108 268 28 280 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=51530 $D=1
M109 269 28 281 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=56160 $D=1
M110 270 28 282 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=60790 $D=1
M111 271 28 283 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=65420 $D=1
M112 8 29 284 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=51530 $D=1
M113 9 29 285 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=56160 $D=1
M114 10 29 286 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=60790 $D=1
M115 11 29 287 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=65420 $D=1
M116 288 30 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=51530 $D=1
M117 289 30 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=56160 $D=1
M118 290 30 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=60790 $D=1
M119 291 30 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=65420 $D=1
M120 292 29 280 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=51530 $D=1
M121 293 29 281 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=56160 $D=1
M122 294 29 282 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=60790 $D=1
M123 295 29 283 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=65420 $D=1
M124 8 292 1234 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=51530 $D=1
M125 9 293 1235 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=56160 $D=1
M126 10 294 1236 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=60790 $D=1
M127 11 295 1237 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=65420 $D=1
M128 296 1234 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=51530 $D=1
M129 297 1235 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=56160 $D=1
M130 298 1236 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=60790 $D=1
M131 299 1237 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=65420 $D=1
M132 292 284 296 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=51530 $D=1
M133 293 285 297 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=56160 $D=1
M134 294 286 298 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=60790 $D=1
M135 295 287 299 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=65420 $D=1
M136 296 30 300 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=51530 $D=1
M137 297 30 301 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=56160 $D=1
M138 298 30 302 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=60790 $D=1
M139 299 30 303 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=65420 $D=1
M140 308 31 296 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=51530 $D=1
M141 309 31 297 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=56160 $D=1
M142 310 31 298 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=60790 $D=1
M143 311 31 299 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=65420 $D=1
M144 304 31 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=51530 $D=1
M145 305 31 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=56160 $D=1
M146 306 31 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=60790 $D=1
M147 307 31 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=65420 $D=1
M148 8 32 312 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=51530 $D=1
M149 9 32 313 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=56160 $D=1
M150 10 32 314 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=60790 $D=1
M151 11 32 315 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=65420 $D=1
M152 316 33 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=51530 $D=1
M153 317 33 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=56160 $D=1
M154 318 33 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=60790 $D=1
M155 319 33 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=65420 $D=1
M156 320 32 280 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=51530 $D=1
M157 321 32 281 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=56160 $D=1
M158 322 32 282 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=60790 $D=1
M159 323 32 283 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=65420 $D=1
M160 8 320 1238 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=51530 $D=1
M161 9 321 1239 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=56160 $D=1
M162 10 322 1240 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=60790 $D=1
M163 11 323 1241 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=65420 $D=1
M164 324 1238 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=51530 $D=1
M165 325 1239 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=56160 $D=1
M166 326 1240 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=60790 $D=1
M167 327 1241 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=65420 $D=1
M168 320 312 324 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=51530 $D=1
M169 321 313 325 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=56160 $D=1
M170 322 314 326 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=60790 $D=1
M171 323 315 327 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=65420 $D=1
M172 324 33 300 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=51530 $D=1
M173 325 33 301 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=56160 $D=1
M174 326 33 302 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=60790 $D=1
M175 327 33 303 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=65420 $D=1
M176 308 34 324 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=51530 $D=1
M177 309 34 325 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=56160 $D=1
M178 310 34 326 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=60790 $D=1
M179 311 34 327 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=65420 $D=1
M180 328 34 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=51530 $D=1
M181 329 34 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=56160 $D=1
M182 330 34 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=60790 $D=1
M183 331 34 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=65420 $D=1
M184 8 35 332 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=51530 $D=1
M185 9 35 333 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=56160 $D=1
M186 10 35 334 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=60790 $D=1
M187 11 35 335 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=65420 $D=1
M188 336 36 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=51530 $D=1
M189 337 36 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=56160 $D=1
M190 338 36 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=60790 $D=1
M191 339 36 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=65420 $D=1
M192 340 35 280 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=51530 $D=1
M193 341 35 281 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=56160 $D=1
M194 342 35 282 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=60790 $D=1
M195 343 35 283 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=65420 $D=1
M196 8 340 1242 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=51530 $D=1
M197 9 341 1243 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=56160 $D=1
M198 10 342 1244 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=60790 $D=1
M199 11 343 1245 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=65420 $D=1
M200 344 1242 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=51530 $D=1
M201 345 1243 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=56160 $D=1
M202 346 1244 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=60790 $D=1
M203 347 1245 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=65420 $D=1
M204 340 332 344 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=51530 $D=1
M205 341 333 345 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=56160 $D=1
M206 342 334 346 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=60790 $D=1
M207 343 335 347 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=65420 $D=1
M208 344 36 300 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=51530 $D=1
M209 345 36 301 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=56160 $D=1
M210 346 36 302 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=60790 $D=1
M211 347 36 303 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=65420 $D=1
M212 308 37 344 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=51530 $D=1
M213 309 37 345 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=56160 $D=1
M214 310 37 346 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=60790 $D=1
M215 311 37 347 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=65420 $D=1
M216 348 37 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=51530 $D=1
M217 349 37 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=56160 $D=1
M218 350 37 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=60790 $D=1
M219 351 37 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=65420 $D=1
M220 8 38 352 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=51530 $D=1
M221 9 38 353 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=56160 $D=1
M222 10 38 354 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=60790 $D=1
M223 11 38 355 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=65420 $D=1
M224 356 39 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=51530 $D=1
M225 357 39 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=56160 $D=1
M226 358 39 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=60790 $D=1
M227 359 39 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=65420 $D=1
M228 360 38 280 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=51530 $D=1
M229 361 38 281 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=56160 $D=1
M230 362 38 282 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=60790 $D=1
M231 363 38 283 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=65420 $D=1
M232 8 360 1246 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=51530 $D=1
M233 9 361 1247 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=56160 $D=1
M234 10 362 1248 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=60790 $D=1
M235 11 363 1249 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=65420 $D=1
M236 364 1246 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=51530 $D=1
M237 365 1247 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=56160 $D=1
M238 366 1248 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=60790 $D=1
M239 367 1249 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=65420 $D=1
M240 360 352 364 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=51530 $D=1
M241 361 353 365 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=56160 $D=1
M242 362 354 366 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=60790 $D=1
M243 363 355 367 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=65420 $D=1
M244 364 39 300 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=51530 $D=1
M245 365 39 301 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=56160 $D=1
M246 366 39 302 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=60790 $D=1
M247 367 39 303 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=65420 $D=1
M248 308 40 364 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=51530 $D=1
M249 309 40 365 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=56160 $D=1
M250 310 40 366 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=60790 $D=1
M251 311 40 367 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=65420 $D=1
M252 368 40 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=51530 $D=1
M253 369 40 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=56160 $D=1
M254 370 40 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=60790 $D=1
M255 371 40 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=65420 $D=1
M256 8 41 372 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=51530 $D=1
M257 9 41 373 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=56160 $D=1
M258 10 41 374 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=60790 $D=1
M259 11 41 375 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=65420 $D=1
M260 376 42 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=51530 $D=1
M261 377 42 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=56160 $D=1
M262 378 42 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=60790 $D=1
M263 379 42 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=65420 $D=1
M264 380 41 280 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=51530 $D=1
M265 381 41 281 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=56160 $D=1
M266 382 41 282 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=60790 $D=1
M267 383 41 283 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=65420 $D=1
M268 8 380 1250 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=51530 $D=1
M269 9 381 1251 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=56160 $D=1
M270 10 382 1252 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=60790 $D=1
M271 11 383 1253 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=65420 $D=1
M272 384 1250 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=51530 $D=1
M273 385 1251 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=56160 $D=1
M274 386 1252 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=60790 $D=1
M275 387 1253 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=65420 $D=1
M276 380 372 384 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=51530 $D=1
M277 381 373 385 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=56160 $D=1
M278 382 374 386 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=60790 $D=1
M279 383 375 387 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=65420 $D=1
M280 384 42 300 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=51530 $D=1
M281 385 42 301 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=56160 $D=1
M282 386 42 302 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=60790 $D=1
M283 387 42 303 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=65420 $D=1
M284 308 43 384 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=51530 $D=1
M285 309 43 385 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=56160 $D=1
M286 310 43 386 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=60790 $D=1
M287 311 43 387 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=65420 $D=1
M288 388 43 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=51530 $D=1
M289 389 43 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=56160 $D=1
M290 390 43 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=60790 $D=1
M291 391 43 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=65420 $D=1
M292 8 44 392 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=51530 $D=1
M293 9 44 393 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=56160 $D=1
M294 10 44 394 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=60790 $D=1
M295 11 44 395 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=65420 $D=1
M296 396 45 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=51530 $D=1
M297 397 45 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=56160 $D=1
M298 398 45 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=60790 $D=1
M299 399 45 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=65420 $D=1
M300 400 44 280 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=51530 $D=1
M301 401 44 281 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=56160 $D=1
M302 402 44 282 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=60790 $D=1
M303 403 44 283 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=65420 $D=1
M304 8 400 1254 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=51530 $D=1
M305 9 401 1255 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=56160 $D=1
M306 10 402 1256 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=60790 $D=1
M307 11 403 1257 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=65420 $D=1
M308 404 1254 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=51530 $D=1
M309 405 1255 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=56160 $D=1
M310 406 1256 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=60790 $D=1
M311 407 1257 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=65420 $D=1
M312 400 392 404 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=51530 $D=1
M313 401 393 405 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=56160 $D=1
M314 402 394 406 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=60790 $D=1
M315 403 395 407 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=65420 $D=1
M316 404 45 300 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=51530 $D=1
M317 405 45 301 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=56160 $D=1
M318 406 45 302 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=60790 $D=1
M319 407 45 303 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=65420 $D=1
M320 308 46 404 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=51530 $D=1
M321 309 46 405 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=56160 $D=1
M322 310 46 406 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=60790 $D=1
M323 311 46 407 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=65420 $D=1
M324 408 46 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=51530 $D=1
M325 409 46 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=56160 $D=1
M326 410 46 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=60790 $D=1
M327 411 46 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=65420 $D=1
M328 8 47 412 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=51530 $D=1
M329 9 47 413 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=56160 $D=1
M330 10 47 414 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=60790 $D=1
M331 11 47 415 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=65420 $D=1
M332 416 48 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=51530 $D=1
M333 417 48 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=56160 $D=1
M334 418 48 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=60790 $D=1
M335 419 48 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=65420 $D=1
M336 420 47 280 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=51530 $D=1
M337 421 47 281 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=56160 $D=1
M338 422 47 282 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=60790 $D=1
M339 423 47 283 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=65420 $D=1
M340 8 420 1258 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=51530 $D=1
M341 9 421 1259 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=56160 $D=1
M342 10 422 1260 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=60790 $D=1
M343 11 423 1261 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=65420 $D=1
M344 424 1258 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=51530 $D=1
M345 425 1259 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=56160 $D=1
M346 426 1260 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=60790 $D=1
M347 427 1261 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=65420 $D=1
M348 420 412 424 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=51530 $D=1
M349 421 413 425 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=56160 $D=1
M350 422 414 426 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=60790 $D=1
M351 423 415 427 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=65420 $D=1
M352 424 48 300 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=51530 $D=1
M353 425 48 301 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=56160 $D=1
M354 426 48 302 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=60790 $D=1
M355 427 48 303 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=65420 $D=1
M356 308 49 424 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=51530 $D=1
M357 309 49 425 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=56160 $D=1
M358 310 49 426 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=60790 $D=1
M359 311 49 427 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=65420 $D=1
M360 428 49 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=51530 $D=1
M361 429 49 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=56160 $D=1
M362 430 49 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=60790 $D=1
M363 431 49 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=65420 $D=1
M364 8 50 432 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=51530 $D=1
M365 9 50 433 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=56160 $D=1
M366 10 50 434 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=60790 $D=1
M367 11 50 435 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=65420 $D=1
M368 436 51 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=51530 $D=1
M369 437 51 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=56160 $D=1
M370 438 51 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=60790 $D=1
M371 439 51 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=65420 $D=1
M372 440 50 280 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=51530 $D=1
M373 441 50 281 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=56160 $D=1
M374 442 50 282 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=60790 $D=1
M375 443 50 283 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=65420 $D=1
M376 8 440 1262 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=51530 $D=1
M377 9 441 1263 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=56160 $D=1
M378 10 442 1264 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=60790 $D=1
M379 11 443 1265 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=65420 $D=1
M380 444 1262 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=51530 $D=1
M381 445 1263 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=56160 $D=1
M382 446 1264 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=60790 $D=1
M383 447 1265 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=65420 $D=1
M384 440 432 444 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=51530 $D=1
M385 441 433 445 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=56160 $D=1
M386 442 434 446 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=60790 $D=1
M387 443 435 447 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=65420 $D=1
M388 444 51 300 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=51530 $D=1
M389 445 51 301 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=56160 $D=1
M390 446 51 302 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=60790 $D=1
M391 447 51 303 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=65420 $D=1
M392 308 52 444 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=51530 $D=1
M393 309 52 445 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=56160 $D=1
M394 310 52 446 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=60790 $D=1
M395 311 52 447 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=65420 $D=1
M396 448 52 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=51530 $D=1
M397 449 52 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=56160 $D=1
M398 450 52 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=60790 $D=1
M399 451 52 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=65420 $D=1
M400 8 53 452 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=51530 $D=1
M401 9 53 453 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=56160 $D=1
M402 10 53 454 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=60790 $D=1
M403 11 53 455 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=65420 $D=1
M404 456 54 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=51530 $D=1
M405 457 54 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=56160 $D=1
M406 458 54 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=60790 $D=1
M407 459 54 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=65420 $D=1
M408 460 53 280 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=51530 $D=1
M409 461 53 281 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=56160 $D=1
M410 462 53 282 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=60790 $D=1
M411 463 53 283 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=65420 $D=1
M412 8 460 1266 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=51530 $D=1
M413 9 461 1267 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=56160 $D=1
M414 10 462 1268 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=60790 $D=1
M415 11 463 1269 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=65420 $D=1
M416 464 1266 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=51530 $D=1
M417 465 1267 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=56160 $D=1
M418 466 1268 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=60790 $D=1
M419 467 1269 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=65420 $D=1
M420 460 452 464 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=51530 $D=1
M421 461 453 465 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=56160 $D=1
M422 462 454 466 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=60790 $D=1
M423 463 455 467 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=65420 $D=1
M424 464 54 300 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=51530 $D=1
M425 465 54 301 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=56160 $D=1
M426 466 54 302 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=60790 $D=1
M427 467 54 303 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=65420 $D=1
M428 308 55 464 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=51530 $D=1
M429 309 55 465 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=56160 $D=1
M430 310 55 466 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=60790 $D=1
M431 311 55 467 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=65420 $D=1
M432 468 55 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=51530 $D=1
M433 469 55 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=56160 $D=1
M434 470 55 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=60790 $D=1
M435 471 55 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=65420 $D=1
M436 8 56 472 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=51530 $D=1
M437 9 56 473 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=56160 $D=1
M438 10 56 474 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=60790 $D=1
M439 11 56 475 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=65420 $D=1
M440 476 57 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=51530 $D=1
M441 477 57 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=56160 $D=1
M442 478 57 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=60790 $D=1
M443 479 57 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=65420 $D=1
M444 480 56 280 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=51530 $D=1
M445 481 56 281 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=56160 $D=1
M446 482 56 282 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=60790 $D=1
M447 483 56 283 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=65420 $D=1
M448 8 480 1270 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=51530 $D=1
M449 9 481 1271 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=56160 $D=1
M450 10 482 1272 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=60790 $D=1
M451 11 483 1273 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=65420 $D=1
M452 484 1270 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=51530 $D=1
M453 485 1271 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=56160 $D=1
M454 486 1272 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=60790 $D=1
M455 487 1273 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=65420 $D=1
M456 480 472 484 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=51530 $D=1
M457 481 473 485 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=56160 $D=1
M458 482 474 486 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=60790 $D=1
M459 483 475 487 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=65420 $D=1
M460 484 57 300 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=51530 $D=1
M461 485 57 301 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=56160 $D=1
M462 486 57 302 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=60790 $D=1
M463 487 57 303 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=65420 $D=1
M464 308 58 484 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=51530 $D=1
M465 309 58 485 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=56160 $D=1
M466 310 58 486 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=60790 $D=1
M467 311 58 487 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=65420 $D=1
M468 488 58 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=51530 $D=1
M469 489 58 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=56160 $D=1
M470 490 58 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=60790 $D=1
M471 491 58 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=65420 $D=1
M472 8 59 492 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=51530 $D=1
M473 9 59 493 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=56160 $D=1
M474 10 59 494 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=60790 $D=1
M475 11 59 495 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=65420 $D=1
M476 496 60 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=51530 $D=1
M477 497 60 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=56160 $D=1
M478 498 60 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=60790 $D=1
M479 499 60 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=65420 $D=1
M480 500 59 280 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=51530 $D=1
M481 501 59 281 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=56160 $D=1
M482 502 59 282 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=60790 $D=1
M483 503 59 283 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=65420 $D=1
M484 8 500 1274 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=51530 $D=1
M485 9 501 1275 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=56160 $D=1
M486 10 502 1276 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=60790 $D=1
M487 11 503 1277 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=65420 $D=1
M488 504 1274 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=51530 $D=1
M489 505 1275 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=56160 $D=1
M490 506 1276 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=60790 $D=1
M491 507 1277 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=65420 $D=1
M492 500 492 504 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=51530 $D=1
M493 501 493 505 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=56160 $D=1
M494 502 494 506 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=60790 $D=1
M495 503 495 507 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=65420 $D=1
M496 504 60 300 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=51530 $D=1
M497 505 60 301 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=56160 $D=1
M498 506 60 302 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=60790 $D=1
M499 507 60 303 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=65420 $D=1
M500 308 61 504 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=51530 $D=1
M501 309 61 505 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=56160 $D=1
M502 310 61 506 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=60790 $D=1
M503 311 61 507 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=65420 $D=1
M504 508 61 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=51530 $D=1
M505 509 61 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=56160 $D=1
M506 510 61 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=60790 $D=1
M507 511 61 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=65420 $D=1
M508 8 62 512 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=51530 $D=1
M509 9 62 513 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=56160 $D=1
M510 10 62 514 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=60790 $D=1
M511 11 62 515 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=65420 $D=1
M512 516 63 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=51530 $D=1
M513 517 63 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=56160 $D=1
M514 518 63 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=60790 $D=1
M515 519 63 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=65420 $D=1
M516 520 62 280 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=51530 $D=1
M517 521 62 281 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=56160 $D=1
M518 522 62 282 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=60790 $D=1
M519 523 62 283 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=65420 $D=1
M520 8 520 1278 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=51530 $D=1
M521 9 521 1279 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=56160 $D=1
M522 10 522 1280 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=60790 $D=1
M523 11 523 1281 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=65420 $D=1
M524 524 1278 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=51530 $D=1
M525 525 1279 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=56160 $D=1
M526 526 1280 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=60790 $D=1
M527 527 1281 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=65420 $D=1
M528 520 512 524 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=51530 $D=1
M529 521 513 525 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=56160 $D=1
M530 522 514 526 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=60790 $D=1
M531 523 515 527 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=65420 $D=1
M532 524 63 300 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=51530 $D=1
M533 525 63 301 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=56160 $D=1
M534 526 63 302 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=60790 $D=1
M535 527 63 303 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=65420 $D=1
M536 308 64 524 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=51530 $D=1
M537 309 64 525 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=56160 $D=1
M538 310 64 526 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=60790 $D=1
M539 311 64 527 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=65420 $D=1
M540 528 64 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=51530 $D=1
M541 529 64 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=56160 $D=1
M542 530 64 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=60790 $D=1
M543 531 64 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=65420 $D=1
M544 8 65 532 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=51530 $D=1
M545 9 65 533 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=56160 $D=1
M546 10 65 534 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=60790 $D=1
M547 11 65 535 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=65420 $D=1
M548 536 66 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=51530 $D=1
M549 537 66 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=56160 $D=1
M550 538 66 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=60790 $D=1
M551 539 66 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=65420 $D=1
M552 540 65 280 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=51530 $D=1
M553 541 65 281 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=56160 $D=1
M554 542 65 282 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=60790 $D=1
M555 543 65 283 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=65420 $D=1
M556 8 540 1282 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=51530 $D=1
M557 9 541 1283 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=56160 $D=1
M558 10 542 1284 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=60790 $D=1
M559 11 543 1285 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=65420 $D=1
M560 544 1282 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=51530 $D=1
M561 545 1283 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=56160 $D=1
M562 546 1284 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=60790 $D=1
M563 547 1285 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=65420 $D=1
M564 540 532 544 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=51530 $D=1
M565 541 533 545 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=56160 $D=1
M566 542 534 546 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=60790 $D=1
M567 543 535 547 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=65420 $D=1
M568 544 66 300 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=51530 $D=1
M569 545 66 301 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=56160 $D=1
M570 546 66 302 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=60790 $D=1
M571 547 66 303 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=65420 $D=1
M572 308 67 544 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=51530 $D=1
M573 309 67 545 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=56160 $D=1
M574 310 67 546 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=60790 $D=1
M575 311 67 547 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=65420 $D=1
M576 548 67 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=51530 $D=1
M577 549 67 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=56160 $D=1
M578 550 67 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=60790 $D=1
M579 551 67 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=65420 $D=1
M580 8 68 552 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=51530 $D=1
M581 9 68 553 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=56160 $D=1
M582 10 68 554 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=60790 $D=1
M583 11 68 555 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=65420 $D=1
M584 556 69 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=51530 $D=1
M585 557 69 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=56160 $D=1
M586 558 69 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=60790 $D=1
M587 559 69 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=65420 $D=1
M588 560 68 280 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=51530 $D=1
M589 561 68 281 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=56160 $D=1
M590 562 68 282 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=60790 $D=1
M591 563 68 283 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=65420 $D=1
M592 8 560 1286 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=51530 $D=1
M593 9 561 1287 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=56160 $D=1
M594 10 562 1288 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=60790 $D=1
M595 11 563 1289 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=65420 $D=1
M596 564 1286 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=51530 $D=1
M597 565 1287 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=56160 $D=1
M598 566 1288 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=60790 $D=1
M599 567 1289 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=65420 $D=1
M600 560 552 564 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=51530 $D=1
M601 561 553 565 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=56160 $D=1
M602 562 554 566 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=60790 $D=1
M603 563 555 567 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=65420 $D=1
M604 564 69 300 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=51530 $D=1
M605 565 69 301 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=56160 $D=1
M606 566 69 302 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=60790 $D=1
M607 567 69 303 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=65420 $D=1
M608 308 70 564 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=51530 $D=1
M609 309 70 565 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=56160 $D=1
M610 310 70 566 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=60790 $D=1
M611 311 70 567 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=65420 $D=1
M612 568 70 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=51530 $D=1
M613 569 70 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=56160 $D=1
M614 570 70 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=60790 $D=1
M615 571 70 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=65420 $D=1
M616 8 71 572 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=51530 $D=1
M617 9 71 573 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=56160 $D=1
M618 10 71 574 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=60790 $D=1
M619 11 71 575 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=65420 $D=1
M620 576 72 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=51530 $D=1
M621 577 72 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=56160 $D=1
M622 578 72 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=60790 $D=1
M623 579 72 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=65420 $D=1
M624 580 71 280 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=51530 $D=1
M625 581 71 281 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=56160 $D=1
M626 582 71 282 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=60790 $D=1
M627 583 71 283 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=65420 $D=1
M628 8 580 1290 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=51530 $D=1
M629 9 581 1291 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=56160 $D=1
M630 10 582 1292 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=60790 $D=1
M631 11 583 1293 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=65420 $D=1
M632 584 1290 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=51530 $D=1
M633 585 1291 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=56160 $D=1
M634 586 1292 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=60790 $D=1
M635 587 1293 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=65420 $D=1
M636 580 572 584 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=51530 $D=1
M637 581 573 585 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=56160 $D=1
M638 582 574 586 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=60790 $D=1
M639 583 575 587 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=65420 $D=1
M640 584 72 300 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=51530 $D=1
M641 585 72 301 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=56160 $D=1
M642 586 72 302 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=60790 $D=1
M643 587 72 303 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=65420 $D=1
M644 308 73 584 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=51530 $D=1
M645 309 73 585 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=56160 $D=1
M646 310 73 586 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=60790 $D=1
M647 311 73 587 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=65420 $D=1
M648 588 73 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=51530 $D=1
M649 589 73 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=56160 $D=1
M650 590 73 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=60790 $D=1
M651 591 73 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=65420 $D=1
M652 8 74 592 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=51530 $D=1
M653 9 74 593 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=56160 $D=1
M654 10 74 594 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=60790 $D=1
M655 11 74 595 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=65420 $D=1
M656 596 75 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=51530 $D=1
M657 597 75 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=56160 $D=1
M658 598 75 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=60790 $D=1
M659 599 75 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=65420 $D=1
M660 600 74 280 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=51530 $D=1
M661 601 74 281 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=56160 $D=1
M662 602 74 282 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=60790 $D=1
M663 603 74 283 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=65420 $D=1
M664 8 600 1294 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=51530 $D=1
M665 9 601 1295 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=56160 $D=1
M666 10 602 1296 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=60790 $D=1
M667 11 603 1297 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=65420 $D=1
M668 604 1294 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=51530 $D=1
M669 605 1295 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=56160 $D=1
M670 606 1296 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=60790 $D=1
M671 607 1297 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=65420 $D=1
M672 600 592 604 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=51530 $D=1
M673 601 593 605 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=56160 $D=1
M674 602 594 606 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=60790 $D=1
M675 603 595 607 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=65420 $D=1
M676 604 75 300 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=51530 $D=1
M677 605 75 301 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=56160 $D=1
M678 606 75 302 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=60790 $D=1
M679 607 75 303 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=65420 $D=1
M680 308 76 604 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=51530 $D=1
M681 309 76 605 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=56160 $D=1
M682 310 76 606 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=60790 $D=1
M683 311 76 607 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=65420 $D=1
M684 608 76 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=51530 $D=1
M685 609 76 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=56160 $D=1
M686 610 76 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=60790 $D=1
M687 611 76 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=65420 $D=1
M688 8 77 612 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=51530 $D=1
M689 9 77 613 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=56160 $D=1
M690 10 77 614 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=60790 $D=1
M691 11 77 615 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=65420 $D=1
M692 616 78 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=51530 $D=1
M693 617 78 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=56160 $D=1
M694 618 78 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=60790 $D=1
M695 619 78 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=65420 $D=1
M696 620 77 280 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=51530 $D=1
M697 621 77 281 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=56160 $D=1
M698 622 77 282 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=60790 $D=1
M699 623 77 283 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=65420 $D=1
M700 8 620 1298 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=51530 $D=1
M701 9 621 1299 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=56160 $D=1
M702 10 622 1300 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=60790 $D=1
M703 11 623 1301 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=65420 $D=1
M704 624 1298 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=51530 $D=1
M705 625 1299 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=56160 $D=1
M706 626 1300 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=60790 $D=1
M707 627 1301 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=65420 $D=1
M708 620 612 624 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=51530 $D=1
M709 621 613 625 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=56160 $D=1
M710 622 614 626 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=60790 $D=1
M711 623 615 627 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=65420 $D=1
M712 624 78 300 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=51530 $D=1
M713 625 78 301 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=56160 $D=1
M714 626 78 302 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=60790 $D=1
M715 627 78 303 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=65420 $D=1
M716 308 79 624 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=51530 $D=1
M717 309 79 625 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=56160 $D=1
M718 310 79 626 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=60790 $D=1
M719 311 79 627 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=65420 $D=1
M720 628 79 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=51530 $D=1
M721 629 79 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=56160 $D=1
M722 630 79 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=60790 $D=1
M723 631 79 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=65420 $D=1
M724 8 80 632 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=51530 $D=1
M725 9 80 633 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=56160 $D=1
M726 10 80 634 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=60790 $D=1
M727 11 80 635 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=65420 $D=1
M728 636 81 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=51530 $D=1
M729 637 81 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=56160 $D=1
M730 638 81 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=60790 $D=1
M731 639 81 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=65420 $D=1
M732 640 80 280 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=51530 $D=1
M733 641 80 281 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=56160 $D=1
M734 642 80 282 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=60790 $D=1
M735 643 80 283 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=65420 $D=1
M736 8 640 1302 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=51530 $D=1
M737 9 641 1303 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=56160 $D=1
M738 10 642 1304 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=60790 $D=1
M739 11 643 1305 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=65420 $D=1
M740 644 1302 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=51530 $D=1
M741 645 1303 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=56160 $D=1
M742 646 1304 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=60790 $D=1
M743 647 1305 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=65420 $D=1
M744 640 632 644 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=51530 $D=1
M745 641 633 645 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=56160 $D=1
M746 642 634 646 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=60790 $D=1
M747 643 635 647 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=65420 $D=1
M748 644 81 300 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=51530 $D=1
M749 645 81 301 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=56160 $D=1
M750 646 81 302 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=60790 $D=1
M751 647 81 303 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=65420 $D=1
M752 308 82 644 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=51530 $D=1
M753 309 82 645 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=56160 $D=1
M754 310 82 646 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=60790 $D=1
M755 311 82 647 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=65420 $D=1
M756 648 82 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=51530 $D=1
M757 649 82 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=56160 $D=1
M758 650 82 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=60790 $D=1
M759 651 82 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=65420 $D=1
M760 8 83 652 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=51530 $D=1
M761 9 83 653 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=56160 $D=1
M762 10 83 654 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=60790 $D=1
M763 11 83 655 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=65420 $D=1
M764 656 84 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=51530 $D=1
M765 657 84 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=56160 $D=1
M766 658 84 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=60790 $D=1
M767 659 84 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=65420 $D=1
M768 660 83 280 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=51530 $D=1
M769 661 83 281 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=56160 $D=1
M770 662 83 282 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=60790 $D=1
M771 663 83 283 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=65420 $D=1
M772 8 660 1306 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=51530 $D=1
M773 9 661 1307 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=56160 $D=1
M774 10 662 1308 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=60790 $D=1
M775 11 663 1309 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=65420 $D=1
M776 664 1306 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=51530 $D=1
M777 665 1307 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=56160 $D=1
M778 666 1308 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=60790 $D=1
M779 667 1309 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=65420 $D=1
M780 660 652 664 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=51530 $D=1
M781 661 653 665 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=56160 $D=1
M782 662 654 666 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=60790 $D=1
M783 663 655 667 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=65420 $D=1
M784 664 84 300 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=51530 $D=1
M785 665 84 301 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=56160 $D=1
M786 666 84 302 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=60790 $D=1
M787 667 84 303 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=65420 $D=1
M788 308 85 664 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=51530 $D=1
M789 309 85 665 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=56160 $D=1
M790 310 85 666 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=60790 $D=1
M791 311 85 667 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=65420 $D=1
M792 668 85 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=51530 $D=1
M793 669 85 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=56160 $D=1
M794 670 85 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=60790 $D=1
M795 671 85 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=65420 $D=1
M796 8 86 672 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=51530 $D=1
M797 9 86 673 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=56160 $D=1
M798 10 86 674 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=60790 $D=1
M799 11 86 675 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=65420 $D=1
M800 676 87 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=51530 $D=1
M801 677 87 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=56160 $D=1
M802 678 87 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=60790 $D=1
M803 679 87 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=65420 $D=1
M804 680 86 280 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=51530 $D=1
M805 681 86 281 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=56160 $D=1
M806 682 86 282 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=60790 $D=1
M807 683 86 283 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=65420 $D=1
M808 8 680 1310 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=51530 $D=1
M809 9 681 1311 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=56160 $D=1
M810 10 682 1312 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=60790 $D=1
M811 11 683 1313 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=65420 $D=1
M812 684 1310 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=51530 $D=1
M813 685 1311 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=56160 $D=1
M814 686 1312 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=60790 $D=1
M815 687 1313 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=65420 $D=1
M816 680 672 684 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=51530 $D=1
M817 681 673 685 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=56160 $D=1
M818 682 674 686 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=60790 $D=1
M819 683 675 687 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=65420 $D=1
M820 684 87 300 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=51530 $D=1
M821 685 87 301 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=56160 $D=1
M822 686 87 302 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=60790 $D=1
M823 687 87 303 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=65420 $D=1
M824 308 88 684 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=51530 $D=1
M825 309 88 685 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=56160 $D=1
M826 310 88 686 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=60790 $D=1
M827 311 88 687 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=65420 $D=1
M828 688 88 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=51530 $D=1
M829 689 88 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=56160 $D=1
M830 690 88 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=60790 $D=1
M831 691 88 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=65420 $D=1
M832 8 89 692 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=51530 $D=1
M833 9 89 693 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=56160 $D=1
M834 10 89 694 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=60790 $D=1
M835 11 89 695 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=65420 $D=1
M836 696 90 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=51530 $D=1
M837 697 90 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=56160 $D=1
M838 698 90 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=60790 $D=1
M839 699 90 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=65420 $D=1
M840 700 89 280 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=51530 $D=1
M841 701 89 281 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=56160 $D=1
M842 702 89 282 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=60790 $D=1
M843 703 89 283 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=65420 $D=1
M844 8 700 1314 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=51530 $D=1
M845 9 701 1315 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=56160 $D=1
M846 10 702 1316 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=60790 $D=1
M847 11 703 1317 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=65420 $D=1
M848 704 1314 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=51530 $D=1
M849 705 1315 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=56160 $D=1
M850 706 1316 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=60790 $D=1
M851 707 1317 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=65420 $D=1
M852 700 692 704 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=51530 $D=1
M853 701 693 705 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=56160 $D=1
M854 702 694 706 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=60790 $D=1
M855 703 695 707 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=65420 $D=1
M856 704 90 300 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=51530 $D=1
M857 705 90 301 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=56160 $D=1
M858 706 90 302 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=60790 $D=1
M859 707 90 303 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=65420 $D=1
M860 308 91 704 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=51530 $D=1
M861 309 91 705 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=56160 $D=1
M862 310 91 706 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=60790 $D=1
M863 311 91 707 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=65420 $D=1
M864 708 91 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=51530 $D=1
M865 709 91 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=56160 $D=1
M866 710 91 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=60790 $D=1
M867 711 91 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=65420 $D=1
M868 8 92 712 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=51530 $D=1
M869 9 92 713 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=56160 $D=1
M870 10 92 714 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=60790 $D=1
M871 11 92 715 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=65420 $D=1
M872 716 93 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=51530 $D=1
M873 717 93 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=56160 $D=1
M874 718 93 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=60790 $D=1
M875 719 93 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=65420 $D=1
M876 720 92 280 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=51530 $D=1
M877 721 92 281 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=56160 $D=1
M878 722 92 282 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=60790 $D=1
M879 723 92 283 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=65420 $D=1
M880 8 720 1318 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=51530 $D=1
M881 9 721 1319 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=56160 $D=1
M882 10 722 1320 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=60790 $D=1
M883 11 723 1321 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=65420 $D=1
M884 724 1318 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=51530 $D=1
M885 725 1319 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=56160 $D=1
M886 726 1320 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=60790 $D=1
M887 727 1321 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=65420 $D=1
M888 720 712 724 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=51530 $D=1
M889 721 713 725 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=56160 $D=1
M890 722 714 726 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=60790 $D=1
M891 723 715 727 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=65420 $D=1
M892 724 93 300 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=51530 $D=1
M893 725 93 301 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=56160 $D=1
M894 726 93 302 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=60790 $D=1
M895 727 93 303 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=65420 $D=1
M896 308 94 724 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=51530 $D=1
M897 309 94 725 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=56160 $D=1
M898 310 94 726 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=60790 $D=1
M899 311 94 727 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=65420 $D=1
M900 728 94 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=51530 $D=1
M901 729 94 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=56160 $D=1
M902 730 94 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=60790 $D=1
M903 731 94 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=65420 $D=1
M904 8 95 732 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=51530 $D=1
M905 9 95 733 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=56160 $D=1
M906 10 95 734 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=60790 $D=1
M907 11 95 735 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=65420 $D=1
M908 736 96 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=51530 $D=1
M909 737 96 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=56160 $D=1
M910 738 96 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=60790 $D=1
M911 739 96 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=65420 $D=1
M912 740 95 280 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=51530 $D=1
M913 741 95 281 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=56160 $D=1
M914 742 95 282 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=60790 $D=1
M915 743 95 283 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=65420 $D=1
M916 8 740 1322 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=51530 $D=1
M917 9 741 1323 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=56160 $D=1
M918 10 742 1324 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=60790 $D=1
M919 11 743 1325 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=65420 $D=1
M920 744 1322 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=51530 $D=1
M921 745 1323 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=56160 $D=1
M922 746 1324 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=60790 $D=1
M923 747 1325 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=65420 $D=1
M924 740 732 744 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=51530 $D=1
M925 741 733 745 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=56160 $D=1
M926 742 734 746 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=60790 $D=1
M927 743 735 747 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=65420 $D=1
M928 744 96 300 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=51530 $D=1
M929 745 96 301 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=56160 $D=1
M930 746 96 302 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=60790 $D=1
M931 747 96 303 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=65420 $D=1
M932 308 97 744 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=51530 $D=1
M933 309 97 745 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=56160 $D=1
M934 310 97 746 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=60790 $D=1
M935 311 97 747 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=65420 $D=1
M936 748 97 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=51530 $D=1
M937 749 97 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=56160 $D=1
M938 750 97 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=60790 $D=1
M939 751 97 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=65420 $D=1
M940 8 98 752 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=51530 $D=1
M941 9 98 753 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=56160 $D=1
M942 10 98 754 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=60790 $D=1
M943 11 98 755 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=65420 $D=1
M944 756 99 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=51530 $D=1
M945 757 99 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=56160 $D=1
M946 758 99 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=60790 $D=1
M947 759 99 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=65420 $D=1
M948 760 98 280 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=51530 $D=1
M949 761 98 281 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=56160 $D=1
M950 762 98 282 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=60790 $D=1
M951 763 98 283 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=65420 $D=1
M952 8 760 1326 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=51530 $D=1
M953 9 761 1327 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=56160 $D=1
M954 10 762 1328 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=60790 $D=1
M955 11 763 1329 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=65420 $D=1
M956 764 1326 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=51530 $D=1
M957 765 1327 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=56160 $D=1
M958 766 1328 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=60790 $D=1
M959 767 1329 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=65420 $D=1
M960 760 752 764 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=51530 $D=1
M961 761 753 765 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=56160 $D=1
M962 762 754 766 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=60790 $D=1
M963 763 755 767 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=65420 $D=1
M964 764 99 300 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=51530 $D=1
M965 765 99 301 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=56160 $D=1
M966 766 99 302 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=60790 $D=1
M967 767 99 303 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=65420 $D=1
M968 308 100 764 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=51530 $D=1
M969 309 100 765 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=56160 $D=1
M970 310 100 766 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=60790 $D=1
M971 311 100 767 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=65420 $D=1
M972 768 100 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=51530 $D=1
M973 769 100 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=56160 $D=1
M974 770 100 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=60790 $D=1
M975 771 100 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=65420 $D=1
M976 8 101 772 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=51530 $D=1
M977 9 101 773 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=56160 $D=1
M978 10 101 774 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=60790 $D=1
M979 11 101 775 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=65420 $D=1
M980 776 102 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=51530 $D=1
M981 777 102 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=56160 $D=1
M982 778 102 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=60790 $D=1
M983 779 102 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=65420 $D=1
M984 780 101 280 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=51530 $D=1
M985 781 101 281 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=56160 $D=1
M986 782 101 282 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=60790 $D=1
M987 783 101 283 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=65420 $D=1
M988 8 780 1330 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=51530 $D=1
M989 9 781 1331 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=56160 $D=1
M990 10 782 1332 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=60790 $D=1
M991 11 783 1333 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=65420 $D=1
M992 784 1330 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=51530 $D=1
M993 785 1331 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=56160 $D=1
M994 786 1332 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=60790 $D=1
M995 787 1333 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=65420 $D=1
M996 780 772 784 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=51530 $D=1
M997 781 773 785 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=56160 $D=1
M998 782 774 786 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=60790 $D=1
M999 783 775 787 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=65420 $D=1
M1000 784 102 300 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=51530 $D=1
M1001 785 102 301 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=56160 $D=1
M1002 786 102 302 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=60790 $D=1
M1003 787 102 303 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=65420 $D=1
M1004 308 103 784 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=51530 $D=1
M1005 309 103 785 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=56160 $D=1
M1006 310 103 786 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=60790 $D=1
M1007 311 103 787 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=65420 $D=1
M1008 788 103 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=51530 $D=1
M1009 789 103 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=56160 $D=1
M1010 790 103 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=60790 $D=1
M1011 791 103 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=65420 $D=1
M1012 8 104 792 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=51530 $D=1
M1013 9 104 793 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=56160 $D=1
M1014 10 104 794 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=60790 $D=1
M1015 11 104 795 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=65420 $D=1
M1016 796 105 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=51530 $D=1
M1017 797 105 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=56160 $D=1
M1018 798 105 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=60790 $D=1
M1019 799 105 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=65420 $D=1
M1020 800 104 280 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=51530 $D=1
M1021 801 104 281 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=56160 $D=1
M1022 802 104 282 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=60790 $D=1
M1023 803 104 283 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=65420 $D=1
M1024 8 800 1334 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=51530 $D=1
M1025 9 801 1335 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=56160 $D=1
M1026 10 802 1336 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=60790 $D=1
M1027 11 803 1337 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=65420 $D=1
M1028 804 1334 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=51530 $D=1
M1029 805 1335 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=56160 $D=1
M1030 806 1336 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=60790 $D=1
M1031 807 1337 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=65420 $D=1
M1032 800 792 804 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=51530 $D=1
M1033 801 793 805 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=56160 $D=1
M1034 802 794 806 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=60790 $D=1
M1035 803 795 807 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=65420 $D=1
M1036 804 105 300 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=51530 $D=1
M1037 805 105 301 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=56160 $D=1
M1038 806 105 302 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=60790 $D=1
M1039 807 105 303 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=65420 $D=1
M1040 308 106 804 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=51530 $D=1
M1041 309 106 805 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=56160 $D=1
M1042 310 106 806 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=60790 $D=1
M1043 311 106 807 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=65420 $D=1
M1044 808 106 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=51530 $D=1
M1045 809 106 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=56160 $D=1
M1046 810 106 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=60790 $D=1
M1047 811 106 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=65420 $D=1
M1048 8 107 812 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=51530 $D=1
M1049 9 107 813 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=56160 $D=1
M1050 10 107 814 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=60790 $D=1
M1051 11 107 815 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=65420 $D=1
M1052 816 108 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=51530 $D=1
M1053 817 108 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=56160 $D=1
M1054 818 108 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=60790 $D=1
M1055 819 108 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=65420 $D=1
M1056 820 107 280 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=51530 $D=1
M1057 821 107 281 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=56160 $D=1
M1058 822 107 282 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=60790 $D=1
M1059 823 107 283 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=65420 $D=1
M1060 8 820 1338 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=51530 $D=1
M1061 9 821 1339 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=56160 $D=1
M1062 10 822 1340 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=60790 $D=1
M1063 11 823 1341 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=65420 $D=1
M1064 824 1338 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=51530 $D=1
M1065 825 1339 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=56160 $D=1
M1066 826 1340 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=60790 $D=1
M1067 827 1341 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=65420 $D=1
M1068 820 812 824 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=51530 $D=1
M1069 821 813 825 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=56160 $D=1
M1070 822 814 826 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=60790 $D=1
M1071 823 815 827 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=65420 $D=1
M1072 824 108 300 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=51530 $D=1
M1073 825 108 301 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=56160 $D=1
M1074 826 108 302 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=60790 $D=1
M1075 827 108 303 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=65420 $D=1
M1076 308 109 824 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=51530 $D=1
M1077 309 109 825 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=56160 $D=1
M1078 310 109 826 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=60790 $D=1
M1079 311 109 827 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=65420 $D=1
M1080 828 109 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=51530 $D=1
M1081 829 109 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=56160 $D=1
M1082 830 109 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=60790 $D=1
M1083 831 109 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=65420 $D=1
M1084 8 110 832 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=51530 $D=1
M1085 9 110 833 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=56160 $D=1
M1086 10 110 834 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=60790 $D=1
M1087 11 110 835 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=65420 $D=1
M1088 836 111 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=51530 $D=1
M1089 837 111 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=56160 $D=1
M1090 838 111 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=60790 $D=1
M1091 839 111 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=65420 $D=1
M1092 840 110 280 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=51530 $D=1
M1093 841 110 281 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=56160 $D=1
M1094 842 110 282 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=60790 $D=1
M1095 843 110 283 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=65420 $D=1
M1096 8 840 1342 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=51530 $D=1
M1097 9 841 1343 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=56160 $D=1
M1098 10 842 1344 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=60790 $D=1
M1099 11 843 1345 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=65420 $D=1
M1100 844 1342 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=51530 $D=1
M1101 845 1343 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=56160 $D=1
M1102 846 1344 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=60790 $D=1
M1103 847 1345 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=65420 $D=1
M1104 840 832 844 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=51530 $D=1
M1105 841 833 845 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=56160 $D=1
M1106 842 834 846 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=60790 $D=1
M1107 843 835 847 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=65420 $D=1
M1108 844 111 300 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=51530 $D=1
M1109 845 111 301 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=56160 $D=1
M1110 846 111 302 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=60790 $D=1
M1111 847 111 303 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=65420 $D=1
M1112 308 112 844 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=51530 $D=1
M1113 309 112 845 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=56160 $D=1
M1114 310 112 846 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=60790 $D=1
M1115 311 112 847 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=65420 $D=1
M1116 848 112 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=51530 $D=1
M1117 849 112 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=56160 $D=1
M1118 850 112 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=60790 $D=1
M1119 851 112 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=65420 $D=1
M1120 8 113 852 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=51530 $D=1
M1121 9 113 853 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=56160 $D=1
M1122 10 113 854 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=60790 $D=1
M1123 11 113 855 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=65420 $D=1
M1124 856 114 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=51530 $D=1
M1125 857 114 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=56160 $D=1
M1126 858 114 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=60790 $D=1
M1127 859 114 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=65420 $D=1
M1128 860 113 280 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=51530 $D=1
M1129 861 113 281 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=56160 $D=1
M1130 862 113 282 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=60790 $D=1
M1131 863 113 283 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=65420 $D=1
M1132 8 860 1346 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=51530 $D=1
M1133 9 861 1347 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=56160 $D=1
M1134 10 862 1348 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=60790 $D=1
M1135 11 863 1349 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=65420 $D=1
M1136 864 1346 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=51530 $D=1
M1137 865 1347 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=56160 $D=1
M1138 866 1348 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=60790 $D=1
M1139 867 1349 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=65420 $D=1
M1140 860 852 864 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=51530 $D=1
M1141 861 853 865 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=56160 $D=1
M1142 862 854 866 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=60790 $D=1
M1143 863 855 867 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=65420 $D=1
M1144 864 114 300 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=51530 $D=1
M1145 865 114 301 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=56160 $D=1
M1146 866 114 302 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=60790 $D=1
M1147 867 114 303 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=65420 $D=1
M1148 308 115 864 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=51530 $D=1
M1149 309 115 865 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=56160 $D=1
M1150 310 115 866 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=60790 $D=1
M1151 311 115 867 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=65420 $D=1
M1152 868 115 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=51530 $D=1
M1153 869 115 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=56160 $D=1
M1154 870 115 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=60790 $D=1
M1155 871 115 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=65420 $D=1
M1156 8 116 872 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=51530 $D=1
M1157 9 116 873 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=56160 $D=1
M1158 10 116 874 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=60790 $D=1
M1159 11 116 875 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=65420 $D=1
M1160 876 117 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=51530 $D=1
M1161 877 117 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=56160 $D=1
M1162 878 117 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=60790 $D=1
M1163 879 117 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=65420 $D=1
M1164 880 116 280 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=51530 $D=1
M1165 881 116 281 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=56160 $D=1
M1166 882 116 282 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=60790 $D=1
M1167 883 116 283 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=65420 $D=1
M1168 8 880 1350 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=51530 $D=1
M1169 9 881 1351 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=56160 $D=1
M1170 10 882 1352 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=60790 $D=1
M1171 11 883 1353 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=65420 $D=1
M1172 884 1350 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=51530 $D=1
M1173 885 1351 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=56160 $D=1
M1174 886 1352 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=60790 $D=1
M1175 887 1353 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=65420 $D=1
M1176 880 872 884 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=51530 $D=1
M1177 881 873 885 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=56160 $D=1
M1178 882 874 886 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=60790 $D=1
M1179 883 875 887 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=65420 $D=1
M1180 884 117 300 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=51530 $D=1
M1181 885 117 301 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=56160 $D=1
M1182 886 117 302 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=60790 $D=1
M1183 887 117 303 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=65420 $D=1
M1184 308 118 884 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=51530 $D=1
M1185 309 118 885 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=56160 $D=1
M1186 310 118 886 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=60790 $D=1
M1187 311 118 887 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=65420 $D=1
M1188 888 118 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=51530 $D=1
M1189 889 118 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=56160 $D=1
M1190 890 118 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=60790 $D=1
M1191 891 118 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=65420 $D=1
M1192 8 119 892 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=51530 $D=1
M1193 9 119 893 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=56160 $D=1
M1194 10 119 894 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=60790 $D=1
M1195 11 119 895 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=65420 $D=1
M1196 896 120 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=51530 $D=1
M1197 897 120 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=56160 $D=1
M1198 898 120 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=60790 $D=1
M1199 899 120 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=65420 $D=1
M1200 900 119 280 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=51530 $D=1
M1201 901 119 281 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=56160 $D=1
M1202 902 119 282 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=60790 $D=1
M1203 903 119 283 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=65420 $D=1
M1204 8 900 1354 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=51530 $D=1
M1205 9 901 1355 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=56160 $D=1
M1206 10 902 1356 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=60790 $D=1
M1207 11 903 1357 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=65420 $D=1
M1208 904 1354 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=51530 $D=1
M1209 905 1355 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=56160 $D=1
M1210 906 1356 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=60790 $D=1
M1211 907 1357 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=65420 $D=1
M1212 900 892 904 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=51530 $D=1
M1213 901 893 905 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=56160 $D=1
M1214 902 894 906 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=60790 $D=1
M1215 903 895 907 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=65420 $D=1
M1216 904 120 300 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=51530 $D=1
M1217 905 120 301 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=56160 $D=1
M1218 906 120 302 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=60790 $D=1
M1219 907 120 303 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=65420 $D=1
M1220 308 121 904 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=51530 $D=1
M1221 309 121 905 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=56160 $D=1
M1222 310 121 906 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=60790 $D=1
M1223 311 121 907 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=65420 $D=1
M1224 908 121 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=51530 $D=1
M1225 909 121 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=56160 $D=1
M1226 910 121 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=60790 $D=1
M1227 911 121 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=65420 $D=1
M1228 8 122 912 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=51530 $D=1
M1229 9 122 913 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=56160 $D=1
M1230 10 122 914 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=60790 $D=1
M1231 11 122 915 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=65420 $D=1
M1232 916 123 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=51530 $D=1
M1233 917 123 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=56160 $D=1
M1234 918 123 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=60790 $D=1
M1235 919 123 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=65420 $D=1
M1236 8 123 300 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=51530 $D=1
M1237 9 123 301 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=56160 $D=1
M1238 10 123 302 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=60790 $D=1
M1239 11 123 303 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=65420 $D=1
M1240 308 122 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=51530 $D=1
M1241 309 122 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=56160 $D=1
M1242 310 122 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=60790 $D=1
M1243 311 122 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=65420 $D=1
M1244 8 924 920 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=51530 $D=1
M1245 9 925 921 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=56160 $D=1
M1246 10 926 922 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=60790 $D=1
M1247 11 927 923 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=65420 $D=1
M1248 924 124 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=51530 $D=1
M1249 925 124 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=56160 $D=1
M1250 926 124 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=60790 $D=1
M1251 927 124 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=65420 $D=1
M1252 1358 300 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=51530 $D=1
M1253 1359 301 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=56160 $D=1
M1254 1360 302 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=60790 $D=1
M1255 1361 303 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=65420 $D=1
M1256 928 920 1358 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=51530 $D=1
M1257 929 921 1359 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=56160 $D=1
M1258 930 922 1360 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=60790 $D=1
M1259 931 923 1361 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=65420 $D=1
M1260 8 928 932 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=51530 $D=1
M1261 9 929 933 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=56160 $D=1
M1262 10 930 934 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=60790 $D=1
M1263 11 931 935 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=65420 $D=1
M1264 1362 932 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=51530 $D=1
M1265 1363 933 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=56160 $D=1
M1266 1364 934 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=60790 $D=1
M1267 1365 935 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=65420 $D=1
M1268 928 924 1362 8 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=51530 $D=1
M1269 929 925 1363 9 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=56160 $D=1
M1270 930 926 1364 10 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=60790 $D=1
M1271 931 927 1365 11 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=65420 $D=1
M1272 8 940 936 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=51530 $D=1
M1273 9 941 937 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=56160 $D=1
M1274 10 942 938 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=60790 $D=1
M1275 11 943 939 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=65420 $D=1
M1276 940 124 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=51530 $D=1
M1277 941 124 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=56160 $D=1
M1278 942 124 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=60790 $D=1
M1279 943 124 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=65420 $D=1
M1280 1366 308 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=51530 $D=1
M1281 1367 309 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=56160 $D=1
M1282 1368 310 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=60790 $D=1
M1283 1369 311 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=65420 $D=1
M1284 944 936 1366 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=51530 $D=1
M1285 945 937 1367 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=56160 $D=1
M1286 946 938 1368 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=60790 $D=1
M1287 947 939 1369 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=65420 $D=1
M1288 8 944 125 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=51530 $D=1
M1289 9 945 126 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=56160 $D=1
M1290 10 946 127 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=60790 $D=1
M1291 11 947 128 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=65420 $D=1
M1292 1370 125 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=51530 $D=1
M1293 1371 126 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=56160 $D=1
M1294 1372 127 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=60790 $D=1
M1295 1373 128 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=65420 $D=1
M1296 944 940 1370 8 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=51530 $D=1
M1297 945 941 1371 9 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=56160 $D=1
M1298 946 942 1372 10 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=60790 $D=1
M1299 947 943 1373 11 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=65420 $D=1
M1300 948 129 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=51530 $D=1
M1301 949 129 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=56160 $D=1
M1302 950 129 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=60790 $D=1
M1303 951 129 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=65420 $D=1
M1304 952 948 932 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=51530 $D=1
M1305 953 949 933 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=56160 $D=1
M1306 954 950 934 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=60790 $D=1
M1307 955 951 935 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=65420 $D=1
M1308 130 129 952 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=51530 $D=1
M1309 131 129 953 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=56160 $D=1
M1310 132 129 954 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=60790 $D=1
M1311 133 129 955 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=65420 $D=1
M1312 956 134 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=51530 $D=1
M1313 957 134 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=56160 $D=1
M1314 958 134 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=60790 $D=1
M1315 959 134 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=65420 $D=1
M1316 960 956 125 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=51530 $D=1
M1317 961 957 126 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=56160 $D=1
M1318 962 958 127 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=60790 $D=1
M1319 963 959 128 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=65420 $D=1
M1320 1374 134 960 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=51530 $D=1
M1321 1375 134 961 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=56160 $D=1
M1322 1376 134 962 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=60790 $D=1
M1323 1377 134 963 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=65420 $D=1
M1324 8 125 1374 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=51530 $D=1
M1325 9 126 1375 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=56160 $D=1
M1326 10 127 1376 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=60790 $D=1
M1327 11 128 1377 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=65420 $D=1
M1328 964 135 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=51530 $D=1
M1329 965 135 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=56160 $D=1
M1330 966 135 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=60790 $D=1
M1331 967 135 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=65420 $D=1
M1332 968 964 960 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=51530 $D=1
M1333 969 965 961 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=56160 $D=1
M1334 970 966 962 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=60790 $D=1
M1335 971 967 963 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=65420 $D=1
M1336 15 135 968 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=51530 $D=1
M1337 16 135 969 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=56160 $D=1
M1338 17 135 970 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=60790 $D=1
M1339 18 135 971 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=65420 $D=1
M1340 975 972 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=51530 $D=1
M1341 976 973 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=56160 $D=1
M1342 977 974 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=60790 $D=1
M1343 978 136 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=65420 $D=1
M1344 8 983 979 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=51530 $D=1
M1345 9 984 980 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=56160 $D=1
M1346 10 985 981 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=60790 $D=1
M1347 11 986 982 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=65420 $D=1
M1348 987 952 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=51530 $D=1
M1349 988 953 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=56160 $D=1
M1350 989 954 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=60790 $D=1
M1351 990 955 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=65420 $D=1
M1352 983 987 972 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=51530 $D=1
M1353 984 988 973 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=56160 $D=1
M1354 985 989 974 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=60790 $D=1
M1355 986 990 136 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=65420 $D=1
M1356 975 952 983 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=51530 $D=1
M1357 976 953 984 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=56160 $D=1
M1358 977 954 985 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=60790 $D=1
M1359 978 955 986 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=65420 $D=1
M1360 991 979 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=51530 $D=1
M1361 992 980 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=56160 $D=1
M1362 993 981 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=60790 $D=1
M1363 994 982 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=65420 $D=1
M1364 137 991 968 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=51530 $D=1
M1365 972 992 969 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=56160 $D=1
M1366 973 993 970 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=60790 $D=1
M1367 974 994 971 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=65420 $D=1
M1368 952 979 137 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=51530 $D=1
M1369 953 980 972 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=56160 $D=1
M1370 954 981 973 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=60790 $D=1
M1371 955 982 974 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=65420 $D=1
M1372 995 137 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=51530 $D=1
M1373 996 972 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=56160 $D=1
M1374 997 973 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=60790 $D=1
M1375 998 974 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=65420 $D=1
M1376 999 979 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=51530 $D=1
M1377 1000 980 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=56160 $D=1
M1378 1001 981 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=60790 $D=1
M1379 1002 982 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=65420 $D=1
M1380 1003 999 995 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=51530 $D=1
M1381 1004 1000 996 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=56160 $D=1
M1382 1005 1001 997 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=60790 $D=1
M1383 1006 1002 998 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=65420 $D=1
M1384 968 979 1003 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=51530 $D=1
M1385 969 980 1004 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=56160 $D=1
M1386 970 981 1005 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=60790 $D=1
M1387 971 982 1006 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=65420 $D=1
M1388 1007 952 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=51530 $D=1
M1389 1008 953 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=56160 $D=1
M1390 1009 954 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=60790 $D=1
M1391 1010 955 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=65420 $D=1
M1392 8 968 1007 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=51530 $D=1
M1393 9 969 1008 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=56160 $D=1
M1394 10 970 1009 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=60790 $D=1
M1395 11 971 1010 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=65420 $D=1
M1396 1011 1003 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=51530 $D=1
M1397 1012 1004 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=56160 $D=1
M1398 1013 1005 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=60790 $D=1
M1399 1014 1006 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=65420 $D=1
M1400 1426 952 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=51530 $D=1
M1401 1427 953 9 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=56160 $D=1
M1402 1428 954 10 10 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=60790 $D=1
M1403 1429 955 11 11 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=65420 $D=1
M1404 1015 968 1426 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=51530 $D=1
M1405 1016 969 1427 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=56160 $D=1
M1406 1017 970 1428 10 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=60790 $D=1
M1407 1018 971 1429 11 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=65420 $D=1
M1408 1430 952 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=51530 $D=1
M1409 1431 953 9 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=56160 $D=1
M1410 1432 954 10 10 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=60790 $D=1
M1411 1433 955 11 11 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=65420 $D=1
M1412 1019 968 1430 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=51530 $D=1
M1413 1020 969 1431 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=56160 $D=1
M1414 1021 970 1432 10 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=60790 $D=1
M1415 1022 971 1433 11 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=65420 $D=1
M1416 1027 952 1023 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=51530 $D=1
M1417 1028 953 1024 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=56160 $D=1
M1418 1029 954 1025 10 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=60790 $D=1
M1419 1030 955 1026 11 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=65420 $D=1
M1420 1023 968 1027 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=51530 $D=1
M1421 1024 969 1028 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=56160 $D=1
M1422 1025 970 1029 10 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=60790 $D=1
M1423 1026 971 1030 11 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=65420 $D=1
M1424 8 1019 1023 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=51530 $D=1
M1425 9 1020 1024 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=56160 $D=1
M1426 10 1021 1025 10 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=60790 $D=1
M1427 11 1022 1026 11 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=65420 $D=1
M1428 1031 144 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=51530 $D=1
M1429 1032 144 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=56160 $D=1
M1430 1033 144 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=60790 $D=1
M1431 1034 144 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=65420 $D=1
M1432 1035 1031 1007 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=51530 $D=1
M1433 1036 1032 1008 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=56160 $D=1
M1434 1037 1033 1009 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=60790 $D=1
M1435 1038 1034 1010 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=65420 $D=1
M1436 1015 144 1035 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=51530 $D=1
M1437 1016 144 1036 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=56160 $D=1
M1438 1017 144 1037 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=60790 $D=1
M1439 1018 144 1038 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=65420 $D=1
M1440 1039 1031 1011 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=51530 $D=1
M1441 1040 1032 1012 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=56160 $D=1
M1442 1041 1033 1013 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=60790 $D=1
M1443 1042 1034 1014 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=65420 $D=1
M1444 1027 144 1039 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=51530 $D=1
M1445 1028 144 1040 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=56160 $D=1
M1446 1029 144 1041 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=60790 $D=1
M1447 1030 144 1042 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=65420 $D=1
M1448 1043 145 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=51530 $D=1
M1449 1044 145 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=56160 $D=1
M1450 1045 145 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=60790 $D=1
M1451 1046 145 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=65420 $D=1
M1452 1047 1043 1039 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=51530 $D=1
M1453 1048 1044 1040 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=56160 $D=1
M1454 1049 1045 1041 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=60790 $D=1
M1455 1050 1046 1042 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=65420 $D=1
M1456 1035 145 1047 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=51530 $D=1
M1457 1036 145 1048 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=56160 $D=1
M1458 1037 145 1049 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=60790 $D=1
M1459 1038 145 1050 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=65420 $D=1
M1460 19 1047 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=51530 $D=1
M1461 20 1048 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=56160 $D=1
M1462 21 1049 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=60790 $D=1
M1463 22 1050 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=65420 $D=1
M1464 1051 146 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=51530 $D=1
M1465 1052 146 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=56160 $D=1
M1466 1053 146 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=60790 $D=1
M1467 1054 146 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=65420 $D=1
M1468 1055 1051 147 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=51530 $D=1
M1469 1056 1052 148 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=56160 $D=1
M1470 1057 1053 149 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=60790 $D=1
M1471 1058 1054 150 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=65420 $D=1
M1472 151 146 1055 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=51530 $D=1
M1473 152 146 1056 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=56160 $D=1
M1474 147 146 1057 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=60790 $D=1
M1475 148 146 1058 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=65420 $D=1
M1476 1059 146 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=51530 $D=1
M1477 1060 146 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=56160 $D=1
M1478 1061 146 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=60790 $D=1
M1479 1062 146 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=65420 $D=1
M1480 1064 1059 153 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=51530 $D=1
M1481 1065 1060 155 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=56160 $D=1
M1482 1066 1061 156 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=60790 $D=1
M1483 1067 1062 158 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=65420 $D=1
M1484 159 146 1064 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=51530 $D=1
M1485 154 146 1065 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=56160 $D=1
M1486 160 146 1066 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=60790 $D=1
M1487 157 146 1067 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=65420 $D=1
M1488 1068 146 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=51530 $D=1
M1489 1069 146 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=56160 $D=1
M1490 1070 146 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=60790 $D=1
M1491 1071 146 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=65420 $D=1
M1492 1072 1068 138 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=51530 $D=1
M1493 1073 1069 143 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=56160 $D=1
M1494 1074 1070 141 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=60790 $D=1
M1495 1075 1071 161 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=65420 $D=1
M1496 162 146 1072 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=51530 $D=1
M1497 163 146 1073 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=56160 $D=1
M1498 164 146 1074 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=60790 $D=1
M1499 165 146 1075 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=65420 $D=1
M1500 1076 146 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=51530 $D=1
M1501 1077 146 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=56160 $D=1
M1502 1078 146 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=60790 $D=1
M1503 1079 146 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=65420 $D=1
M1504 1080 1076 166 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=51530 $D=1
M1505 1081 1077 167 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=56160 $D=1
M1506 1082 1078 168 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=60790 $D=1
M1507 1083 1079 169 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=65420 $D=1
M1508 170 146 1080 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=51530 $D=1
M1509 171 146 1081 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=56160 $D=1
M1510 172 146 1082 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=60790 $D=1
M1511 173 146 1083 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=65420 $D=1
M1512 1084 146 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=51530 $D=1
M1513 1085 146 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=56160 $D=1
M1514 1086 146 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=60790 $D=1
M1515 1087 146 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=65420 $D=1
M1516 1088 1084 174 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=51530 $D=1
M1517 1089 1085 175 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=56160 $D=1
M1518 1090 1086 176 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=60790 $D=1
M1519 1091 1087 177 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=65420 $D=1
M1520 178 146 1088 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=51530 $D=1
M1521 178 146 1089 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=56160 $D=1
M1522 178 146 1090 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=60790 $D=1
M1523 178 146 1091 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=65420 $D=1
M1524 8 952 1390 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=51530 $D=1
M1525 9 953 1391 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=56160 $D=1
M1526 10 954 1392 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=60790 $D=1
M1527 11 955 1393 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=65420 $D=1
M1528 152 1390 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=51530 $D=1
M1529 147 1391 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=56160 $D=1
M1530 148 1392 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=60790 $D=1
M1531 149 1393 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=65420 $D=1
M1532 1092 179 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=51530 $D=1
M1533 1093 179 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=56160 $D=1
M1534 1094 179 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=60790 $D=1
M1535 1095 179 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=65420 $D=1
M1536 160 1092 152 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=51530 $D=1
M1537 157 1093 147 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=56160 $D=1
M1538 153 1094 148 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=60790 $D=1
M1539 155 1095 149 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=65420 $D=1
M1540 1055 179 160 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=51530 $D=1
M1541 1056 179 157 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=56160 $D=1
M1542 1057 179 153 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=60790 $D=1
M1543 1058 179 155 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=65420 $D=1
M1544 1096 180 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=51530 $D=1
M1545 1097 180 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=56160 $D=1
M1546 1098 180 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=60790 $D=1
M1547 1099 180 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=65420 $D=1
M1548 181 1096 160 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=51530 $D=1
M1549 142 1097 157 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=56160 $D=1
M1550 140 1098 153 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=60790 $D=1
M1551 139 1099 155 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=65420 $D=1
M1552 1064 180 181 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=51530 $D=1
M1553 1065 180 142 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=56160 $D=1
M1554 1066 180 140 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=60790 $D=1
M1555 1067 180 139 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=65420 $D=1
M1556 1100 182 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=51530 $D=1
M1557 1101 182 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=56160 $D=1
M1558 1102 182 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=60790 $D=1
M1559 1103 182 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=65420 $D=1
M1560 183 1100 181 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=51530 $D=1
M1561 184 1101 142 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=56160 $D=1
M1562 185 1102 140 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=60790 $D=1
M1563 186 1103 139 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=65420 $D=1
M1564 1072 182 183 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=51530 $D=1
M1565 1073 182 184 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=56160 $D=1
M1566 1074 182 185 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=60790 $D=1
M1567 1075 182 186 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=65420 $D=1
M1568 1104 187 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=51530 $D=1
M1569 1105 187 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=56160 $D=1
M1570 1106 187 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=60790 $D=1
M1571 1107 187 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=65420 $D=1
M1572 188 1104 183 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=51530 $D=1
M1573 189 1105 184 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=56160 $D=1
M1574 190 1106 185 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=60790 $D=1
M1575 191 1107 186 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=65420 $D=1
M1576 1080 187 188 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=51530 $D=1
M1577 1081 187 189 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=56160 $D=1
M1578 1082 187 190 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=60790 $D=1
M1579 1083 187 191 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=65420 $D=1
M1580 1108 192 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=51530 $D=1
M1581 1109 192 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=56160 $D=1
M1582 1110 192 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=60790 $D=1
M1583 1111 192 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=65420 $D=1
M1584 23 1108 188 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=51530 $D=1
M1585 24 1109 189 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=56160 $D=1
M1586 25 1110 190 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=60790 $D=1
M1587 26 1111 191 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=65420 $D=1
M1588 1088 192 23 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=51530 $D=1
M1589 1089 192 24 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=56160 $D=1
M1590 1090 192 25 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=60790 $D=1
M1591 1091 192 26 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=65420 $D=1
M1592 1112 193 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=51530 $D=1
M1593 1113 193 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=56160 $D=1
M1594 1114 193 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=60790 $D=1
M1595 1115 193 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=65420 $D=1
M1596 1116 1112 125 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=51530 $D=1
M1597 1117 1113 126 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=56160 $D=1
M1598 1118 1114 127 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=60790 $D=1
M1599 1119 1115 128 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=65420 $D=1
M1600 15 193 1116 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=51530 $D=1
M1601 16 193 1117 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=56160 $D=1
M1602 17 193 1118 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=60790 $D=1
M1603 18 193 1119 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=65420 $D=1
M1604 1434 932 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=51530 $D=1
M1605 1435 933 9 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=56160 $D=1
M1606 1436 934 10 10 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=60790 $D=1
M1607 1437 935 11 11 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=65420 $D=1
M1608 1120 1116 1434 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=51530 $D=1
M1609 1121 1117 1435 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=56160 $D=1
M1610 1122 1118 1436 10 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=60790 $D=1
M1611 1123 1119 1437 11 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=65420 $D=1
M1612 1128 932 1124 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=51530 $D=1
M1613 1129 933 1125 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=56160 $D=1
M1614 1130 934 1126 10 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=60790 $D=1
M1615 1131 935 1127 11 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=65420 $D=1
M1616 1124 1116 1128 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=51530 $D=1
M1617 1125 1117 1129 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=56160 $D=1
M1618 1126 1118 1130 10 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=60790 $D=1
M1619 1127 1119 1131 11 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=65420 $D=1
M1620 8 1120 1124 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=51530 $D=1
M1621 9 1121 1125 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=56160 $D=1
M1622 10 1122 1126 10 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=60790 $D=1
M1623 11 1123 1127 11 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=65420 $D=1
M1624 1438 194 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=51530 $D=1
M1625 1439 1132 9 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=56160 $D=1
M1626 1440 1133 10 10 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=60790 $D=1
M1627 1441 1134 11 11 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=65420 $D=1
M1628 1394 1128 1438 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=51530 $D=1
M1629 1395 1129 1439 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=56160 $D=1
M1630 1396 1130 1440 10 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=60790 $D=1
M1631 1397 1131 1441 11 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=65420 $D=1
M1632 1132 1394 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=51530 $D=1
M1633 1135 1395 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=56160 $D=1
M1634 1134 1396 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=60790 $D=1
M1635 195 1397 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=65420 $D=1
M1636 1136 932 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=51530 $D=1
M1637 1137 933 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=56160 $D=1
M1638 1138 934 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=60790 $D=1
M1639 1139 935 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=65420 $D=1
M1640 8 1140 1136 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=51530 $D=1
M1641 9 1141 1137 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=56160 $D=1
M1642 10 1142 1138 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=60790 $D=1
M1643 11 1143 1139 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=65420 $D=1
M1644 1140 1116 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=51530 $D=1
M1645 1141 1117 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=56160 $D=1
M1646 1142 1118 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=60790 $D=1
M1647 1143 1119 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=65420 $D=1
M1648 1442 1136 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=51530 $D=1
M1649 1443 1137 9 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=56160 $D=1
M1650 1444 1138 10 10 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=60790 $D=1
M1651 1445 1139 11 11 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=65420 $D=1
M1652 1144 194 1442 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=51530 $D=1
M1653 1145 1132 1443 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=56160 $D=1
M1654 1146 1133 1444 10 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=60790 $D=1
M1655 1147 1134 1445 11 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=65420 $D=1
M1656 1151 196 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=51530 $D=1
M1657 1152 1148 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=56160 $D=1
M1658 1153 1149 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=60790 $D=1
M1659 1154 1150 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=65420 $D=1
M1660 1446 1144 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=51530 $D=1
M1661 1447 1145 9 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=56160 $D=1
M1662 1448 1146 10 10 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=60790 $D=1
M1663 1449 1147 11 11 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=65420 $D=1
M1664 1148 1151 1446 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=51530 $D=1
M1665 1149 1152 1447 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=56160 $D=1
M1666 1150 1153 1448 10 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=60790 $D=1
M1667 197 1154 1449 11 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=65420 $D=1
M1668 1158 1155 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=51530 $D=1
M1669 1159 1156 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=56160 $D=1
M1670 1160 1157 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=60790 $D=1
M1671 1161 198 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=65420 $D=1
M1672 8 1166 1162 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=51530 $D=1
M1673 9 1167 1163 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=56160 $D=1
M1674 10 1168 1164 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=60790 $D=1
M1675 11 1169 1165 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=65420 $D=1
M1676 1170 130 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=51530 $D=1
M1677 1171 131 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=56160 $D=1
M1678 1172 132 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=60790 $D=1
M1679 1173 133 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=65420 $D=1
M1680 1166 1170 1155 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=51530 $D=1
M1681 1167 1171 1156 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=56160 $D=1
M1682 1168 1172 1157 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=60790 $D=1
M1683 1169 1173 198 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=65420 $D=1
M1684 1158 130 1166 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=51530 $D=1
M1685 1159 131 1167 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=56160 $D=1
M1686 1160 132 1168 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=60790 $D=1
M1687 1161 133 1169 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=65420 $D=1
M1688 1174 1162 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=51530 $D=1
M1689 1175 1163 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=56160 $D=1
M1690 1176 1164 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=60790 $D=1
M1691 1177 1165 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=65420 $D=1
M1692 199 1174 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=51530 $D=1
M1693 1155 1175 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=56160 $D=1
M1694 1156 1176 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=60790 $D=1
M1695 1157 1177 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=65420 $D=1
M1696 130 1162 199 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=51530 $D=1
M1697 131 1163 1155 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=56160 $D=1
M1698 132 1164 1156 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=60790 $D=1
M1699 133 1165 1157 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=65420 $D=1
M1700 1178 199 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=51530 $D=1
M1701 1179 1155 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=56160 $D=1
M1702 1180 1156 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=60790 $D=1
M1703 1181 1157 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=65420 $D=1
M1704 1182 1162 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=51530 $D=1
M1705 1183 1163 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=56160 $D=1
M1706 1184 1164 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=60790 $D=1
M1707 1185 1165 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=65420 $D=1
M1708 256 1182 1178 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=51530 $D=1
M1709 257 1183 1179 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=56160 $D=1
M1710 258 1184 1180 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=60790 $D=1
M1711 259 1185 1181 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=65420 $D=1
M1712 8 1162 256 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=51530 $D=1
M1713 9 1163 257 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=56160 $D=1
M1714 10 1164 258 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=60790 $D=1
M1715 11 1165 259 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=65420 $D=1
M1716 1186 200 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=51530 $D=1
M1717 1187 200 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=56160 $D=1
M1718 1188 200 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=60790 $D=1
M1719 1189 200 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=65420 $D=1
M1720 1190 1186 256 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=51530 $D=1
M1721 1191 1187 257 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=56160 $D=1
M1722 1192 1188 258 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=60790 $D=1
M1723 1193 1189 259 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=65420 $D=1
M1724 19 200 1190 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=51530 $D=1
M1725 20 200 1191 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=56160 $D=1
M1726 21 200 1192 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=60790 $D=1
M1727 22 200 1193 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=65420 $D=1
M1728 1194 201 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=51530 $D=1
M1729 1195 201 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=56160 $D=1
M1730 1196 201 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=60790 $D=1
M1731 1197 201 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=65420 $D=1
M1732 201 1194 1190 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=51530 $D=1
M1733 201 1195 1191 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=56160 $D=1
M1734 201 1196 1192 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=60790 $D=1
M1735 201 1197 1193 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=65420 $D=1
M1736 8 201 201 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=51530 $D=1
M1737 9 201 201 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=56160 $D=1
M1738 10 201 201 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=60790 $D=1
M1739 11 201 201 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=65420 $D=1
M1740 1198 124 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=51530 $D=1
M1741 1199 124 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=56160 $D=1
M1742 1200 124 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=60790 $D=1
M1743 1201 124 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=65420 $D=1
M1744 8 1198 1202 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=51530 $D=1
M1745 9 1199 1203 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=56160 $D=1
M1746 10 1200 1204 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=60790 $D=1
M1747 11 1201 1205 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=65420 $D=1
M1748 1206 124 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=51530 $D=1
M1749 1207 124 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=56160 $D=1
M1750 1208 124 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=60790 $D=1
M1751 1209 124 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=65420 $D=1
M1752 1210 1198 201 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=51530 $D=1
M1753 1211 1199 201 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=56160 $D=1
M1754 1212 1200 201 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=60790 $D=1
M1755 1213 1201 201 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=65420 $D=1
M1756 8 1210 1398 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=51530 $D=1
M1757 9 1211 1399 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=56160 $D=1
M1758 10 1212 1400 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=60790 $D=1
M1759 11 1213 1401 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=65420 $D=1
M1760 1214 1398 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=51530 $D=1
M1761 1215 1399 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=56160 $D=1
M1762 1216 1400 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=60790 $D=1
M1763 1217 1401 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=65420 $D=1
M1764 1210 1202 1214 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=51530 $D=1
M1765 1211 1203 1215 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=56160 $D=1
M1766 1212 1204 1216 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=60790 $D=1
M1767 1213 1205 1217 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=65420 $D=1
M1768 1218 124 1214 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=51530 $D=1
M1769 1219 124 1215 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=56160 $D=1
M1770 1220 124 1216 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=60790 $D=1
M1771 1221 124 1217 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=65420 $D=1
M1772 8 1226 1222 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=51530 $D=1
M1773 9 1227 1223 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=56160 $D=1
M1774 10 1228 1224 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=60790 $D=1
M1775 11 1229 1225 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=65420 $D=1
M1776 1226 124 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=51530 $D=1
M1777 1227 124 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=56160 $D=1
M1778 1228 124 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=60790 $D=1
M1779 1229 124 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=65420 $D=1
M1780 1402 1218 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=51530 $D=1
M1781 1403 1219 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=56160 $D=1
M1782 1404 1220 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=60790 $D=1
M1783 1405 1221 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=65420 $D=1
M1784 1230 1222 1402 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=51530 $D=1
M1785 1231 1223 1403 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=56160 $D=1
M1786 1232 1224 1404 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=60790 $D=1
M1787 1233 1225 1405 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=65420 $D=1
M1788 8 1230 130 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=51530 $D=1
M1789 9 1231 131 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=56160 $D=1
M1790 10 1232 132 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=60790 $D=1
M1791 11 1233 133 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=65420 $D=1
M1792 1406 130 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=51530 $D=1
M1793 1407 131 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=56160 $D=1
M1794 1408 132 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=60790 $D=1
M1795 1409 133 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=65420 $D=1
M1796 1230 1226 1406 8 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=51530 $D=1
M1797 1231 1227 1407 9 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=56160 $D=1
M1798 1232 1228 1408 10 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=60790 $D=1
M1799 1233 1229 1409 11 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=65420 $D=1
M1800 208 1 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=52780 $D=0
M1801 209 1 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=57410 $D=0
M1802 210 1 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=62040 $D=0
M1803 211 1 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=66670 $D=0
M1804 212 1 2 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=52780 $D=0
M1805 213 1 3 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=57410 $D=0
M1806 214 1 4 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=62040 $D=0
M1807 215 1 5 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=66670 $D=0
M1808 8 208 212 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=52780 $D=0
M1809 9 209 213 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=57410 $D=0
M1810 10 210 214 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=62040 $D=0
M1811 11 211 215 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=66670 $D=0
M1812 216 1 6 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=52780 $D=0
M1813 217 1 6 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=57410 $D=0
M1814 218 1 6 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=62040 $D=0
M1815 219 1 6 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=66670 $D=0
M1816 7 208 216 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=52780 $D=0
M1817 7 209 217 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=57410 $D=0
M1818 7 210 218 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=62040 $D=0
M1819 7 211 219 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=66670 $D=0
M1820 220 1 8 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=52780 $D=0
M1821 221 1 9 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=57410 $D=0
M1822 222 1 10 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=62040 $D=0
M1823 223 1 11 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=66670 $D=0
M1824 8 208 220 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=52780 $D=0
M1825 9 209 221 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=57410 $D=0
M1826 10 210 222 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=62040 $D=0
M1827 11 211 223 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=66670 $D=0
M1828 228 12 220 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=52780 $D=0
M1829 229 12 221 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=57410 $D=0
M1830 230 12 222 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=62040 $D=0
M1831 231 12 223 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=66670 $D=0
M1832 224 12 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=52780 $D=0
M1833 225 12 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=57410 $D=0
M1834 226 12 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=62040 $D=0
M1835 227 12 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=66670 $D=0
M1836 232 12 216 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=52780 $D=0
M1837 233 12 217 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=57410 $D=0
M1838 234 12 218 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=62040 $D=0
M1839 235 12 219 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=66670 $D=0
M1840 212 224 232 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=52780 $D=0
M1841 213 225 233 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=57410 $D=0
M1842 214 226 234 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=62040 $D=0
M1843 215 227 235 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=66670 $D=0
M1844 236 13 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=52780 $D=0
M1845 237 13 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=57410 $D=0
M1846 238 13 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=62040 $D=0
M1847 239 13 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=66670 $D=0
M1848 240 13 232 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=52780 $D=0
M1849 241 13 233 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=57410 $D=0
M1850 242 13 234 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=62040 $D=0
M1851 243 13 235 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=66670 $D=0
M1852 228 236 240 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=52780 $D=0
M1853 229 237 241 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=57410 $D=0
M1854 230 238 242 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=62040 $D=0
M1855 231 239 243 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=66670 $D=0
M1856 244 14 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=52780 $D=0
M1857 245 14 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=57410 $D=0
M1858 246 14 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=62040 $D=0
M1859 247 14 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=66670 $D=0
M1860 248 14 8 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=52780 $D=0
M1861 249 14 9 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=57410 $D=0
M1862 250 14 10 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=62040 $D=0
M1863 251 14 11 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=66670 $D=0
M1864 15 244 248 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=52780 $D=0
M1865 16 245 249 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=57410 $D=0
M1866 17 246 250 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=62040 $D=0
M1867 18 247 251 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=66670 $D=0
M1868 252 14 19 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=52780 $D=0
M1869 253 14 20 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=57410 $D=0
M1870 254 14 21 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=62040 $D=0
M1871 255 14 22 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=66670 $D=0
M1872 23 244 252 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=52780 $D=0
M1873 24 245 253 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=57410 $D=0
M1874 25 246 254 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=62040 $D=0
M1875 26 247 255 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=66670 $D=0
M1876 260 14 256 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=52780 $D=0
M1877 261 14 257 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=57410 $D=0
M1878 262 14 258 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=62040 $D=0
M1879 263 14 259 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=66670 $D=0
M1880 240 244 260 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=52780 $D=0
M1881 241 245 261 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=57410 $D=0
M1882 242 246 262 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=62040 $D=0
M1883 243 247 263 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=66670 $D=0
M1884 268 27 260 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=52780 $D=0
M1885 269 27 261 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=57410 $D=0
M1886 270 27 262 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=62040 $D=0
M1887 271 27 263 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=66670 $D=0
M1888 264 27 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=52780 $D=0
M1889 265 27 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=57410 $D=0
M1890 266 27 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=62040 $D=0
M1891 267 27 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=66670 $D=0
M1892 272 27 252 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=52780 $D=0
M1893 273 27 253 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=57410 $D=0
M1894 274 27 254 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=62040 $D=0
M1895 275 27 255 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=66670 $D=0
M1896 248 264 272 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=52780 $D=0
M1897 249 265 273 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=57410 $D=0
M1898 250 266 274 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=62040 $D=0
M1899 251 267 275 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=66670 $D=0
M1900 276 28 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=52780 $D=0
M1901 277 28 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=57410 $D=0
M1902 278 28 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=62040 $D=0
M1903 279 28 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=66670 $D=0
M1904 280 28 272 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=52780 $D=0
M1905 281 28 273 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=57410 $D=0
M1906 282 28 274 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=62040 $D=0
M1907 283 28 275 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=66670 $D=0
M1908 268 276 280 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=52780 $D=0
M1909 269 277 281 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=57410 $D=0
M1910 270 278 282 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=62040 $D=0
M1911 271 279 283 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=66670 $D=0
M1912 202 29 284 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=52780 $D=0
M1913 203 29 285 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=57410 $D=0
M1914 204 29 286 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=62040 $D=0
M1915 205 29 287 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=66670 $D=0
M1916 288 30 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=52780 $D=0
M1917 289 30 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=57410 $D=0
M1918 290 30 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=62040 $D=0
M1919 291 30 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=66670 $D=0
M1920 292 284 280 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=52780 $D=0
M1921 293 285 281 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=57410 $D=0
M1922 294 286 282 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=62040 $D=0
M1923 295 287 283 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=66670 $D=0
M1924 202 292 1234 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=52780 $D=0
M1925 203 293 1235 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=57410 $D=0
M1926 204 294 1236 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=62040 $D=0
M1927 205 295 1237 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=66670 $D=0
M1928 296 1234 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=52780 $D=0
M1929 297 1235 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=57410 $D=0
M1930 298 1236 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=62040 $D=0
M1931 299 1237 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=66670 $D=0
M1932 292 29 296 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=52780 $D=0
M1933 293 29 297 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=57410 $D=0
M1934 294 29 298 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=62040 $D=0
M1935 295 29 299 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=66670 $D=0
M1936 296 288 300 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=52780 $D=0
M1937 297 289 301 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=57410 $D=0
M1938 298 290 302 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=62040 $D=0
M1939 299 291 303 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=66670 $D=0
M1940 308 304 296 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=52780 $D=0
M1941 309 305 297 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=57410 $D=0
M1942 310 306 298 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=62040 $D=0
M1943 311 307 299 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=66670 $D=0
M1944 304 31 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=52780 $D=0
M1945 305 31 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=57410 $D=0
M1946 306 31 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=62040 $D=0
M1947 307 31 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=66670 $D=0
M1948 202 32 312 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=52780 $D=0
M1949 203 32 313 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=57410 $D=0
M1950 204 32 314 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=62040 $D=0
M1951 205 32 315 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=66670 $D=0
M1952 316 33 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=52780 $D=0
M1953 317 33 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=57410 $D=0
M1954 318 33 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=62040 $D=0
M1955 319 33 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=66670 $D=0
M1956 320 312 280 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=52780 $D=0
M1957 321 313 281 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=57410 $D=0
M1958 322 314 282 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=62040 $D=0
M1959 323 315 283 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=66670 $D=0
M1960 202 320 1238 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=52780 $D=0
M1961 203 321 1239 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=57410 $D=0
M1962 204 322 1240 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=62040 $D=0
M1963 205 323 1241 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=66670 $D=0
M1964 324 1238 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=52780 $D=0
M1965 325 1239 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=57410 $D=0
M1966 326 1240 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=62040 $D=0
M1967 327 1241 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=66670 $D=0
M1968 320 32 324 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=52780 $D=0
M1969 321 32 325 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=57410 $D=0
M1970 322 32 326 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=62040 $D=0
M1971 323 32 327 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=66670 $D=0
M1972 324 316 300 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=52780 $D=0
M1973 325 317 301 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=57410 $D=0
M1974 326 318 302 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=62040 $D=0
M1975 327 319 303 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=66670 $D=0
M1976 308 328 324 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=52780 $D=0
M1977 309 329 325 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=57410 $D=0
M1978 310 330 326 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=62040 $D=0
M1979 311 331 327 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=66670 $D=0
M1980 328 34 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=52780 $D=0
M1981 329 34 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=57410 $D=0
M1982 330 34 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=62040 $D=0
M1983 331 34 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=66670 $D=0
M1984 202 35 332 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=52780 $D=0
M1985 203 35 333 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=57410 $D=0
M1986 204 35 334 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=62040 $D=0
M1987 205 35 335 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=66670 $D=0
M1988 336 36 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=52780 $D=0
M1989 337 36 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=57410 $D=0
M1990 338 36 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=62040 $D=0
M1991 339 36 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=66670 $D=0
M1992 340 332 280 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=52780 $D=0
M1993 341 333 281 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=57410 $D=0
M1994 342 334 282 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=62040 $D=0
M1995 343 335 283 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=66670 $D=0
M1996 202 340 1242 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=52780 $D=0
M1997 203 341 1243 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=57410 $D=0
M1998 204 342 1244 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=62040 $D=0
M1999 205 343 1245 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=66670 $D=0
M2000 344 1242 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=52780 $D=0
M2001 345 1243 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=57410 $D=0
M2002 346 1244 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=62040 $D=0
M2003 347 1245 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=66670 $D=0
M2004 340 35 344 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=52780 $D=0
M2005 341 35 345 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=57410 $D=0
M2006 342 35 346 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=62040 $D=0
M2007 343 35 347 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=66670 $D=0
M2008 344 336 300 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=52780 $D=0
M2009 345 337 301 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=57410 $D=0
M2010 346 338 302 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=62040 $D=0
M2011 347 339 303 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=66670 $D=0
M2012 308 348 344 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=52780 $D=0
M2013 309 349 345 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=57410 $D=0
M2014 310 350 346 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=62040 $D=0
M2015 311 351 347 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=66670 $D=0
M2016 348 37 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=52780 $D=0
M2017 349 37 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=57410 $D=0
M2018 350 37 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=62040 $D=0
M2019 351 37 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=66670 $D=0
M2020 202 38 352 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=52780 $D=0
M2021 203 38 353 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=57410 $D=0
M2022 204 38 354 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=62040 $D=0
M2023 205 38 355 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=66670 $D=0
M2024 356 39 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=52780 $D=0
M2025 357 39 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=57410 $D=0
M2026 358 39 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=62040 $D=0
M2027 359 39 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=66670 $D=0
M2028 360 352 280 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=52780 $D=0
M2029 361 353 281 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=57410 $D=0
M2030 362 354 282 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=62040 $D=0
M2031 363 355 283 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=66670 $D=0
M2032 202 360 1246 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=52780 $D=0
M2033 203 361 1247 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=57410 $D=0
M2034 204 362 1248 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=62040 $D=0
M2035 205 363 1249 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=66670 $D=0
M2036 364 1246 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=52780 $D=0
M2037 365 1247 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=57410 $D=0
M2038 366 1248 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=62040 $D=0
M2039 367 1249 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=66670 $D=0
M2040 360 38 364 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=52780 $D=0
M2041 361 38 365 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=57410 $D=0
M2042 362 38 366 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=62040 $D=0
M2043 363 38 367 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=66670 $D=0
M2044 364 356 300 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=52780 $D=0
M2045 365 357 301 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=57410 $D=0
M2046 366 358 302 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=62040 $D=0
M2047 367 359 303 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=66670 $D=0
M2048 308 368 364 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=52780 $D=0
M2049 309 369 365 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=57410 $D=0
M2050 310 370 366 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=62040 $D=0
M2051 311 371 367 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=66670 $D=0
M2052 368 40 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=52780 $D=0
M2053 369 40 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=57410 $D=0
M2054 370 40 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=62040 $D=0
M2055 371 40 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=66670 $D=0
M2056 202 41 372 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=52780 $D=0
M2057 203 41 373 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=57410 $D=0
M2058 204 41 374 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=62040 $D=0
M2059 205 41 375 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=66670 $D=0
M2060 376 42 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=52780 $D=0
M2061 377 42 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=57410 $D=0
M2062 378 42 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=62040 $D=0
M2063 379 42 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=66670 $D=0
M2064 380 372 280 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=52780 $D=0
M2065 381 373 281 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=57410 $D=0
M2066 382 374 282 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=62040 $D=0
M2067 383 375 283 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=66670 $D=0
M2068 202 380 1250 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=52780 $D=0
M2069 203 381 1251 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=57410 $D=0
M2070 204 382 1252 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=62040 $D=0
M2071 205 383 1253 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=66670 $D=0
M2072 384 1250 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=52780 $D=0
M2073 385 1251 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=57410 $D=0
M2074 386 1252 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=62040 $D=0
M2075 387 1253 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=66670 $D=0
M2076 380 41 384 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=52780 $D=0
M2077 381 41 385 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=57410 $D=0
M2078 382 41 386 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=62040 $D=0
M2079 383 41 387 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=66670 $D=0
M2080 384 376 300 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=52780 $D=0
M2081 385 377 301 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=57410 $D=0
M2082 386 378 302 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=62040 $D=0
M2083 387 379 303 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=66670 $D=0
M2084 308 388 384 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=52780 $D=0
M2085 309 389 385 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=57410 $D=0
M2086 310 390 386 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=62040 $D=0
M2087 311 391 387 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=66670 $D=0
M2088 388 43 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=52780 $D=0
M2089 389 43 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=57410 $D=0
M2090 390 43 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=62040 $D=0
M2091 391 43 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=66670 $D=0
M2092 202 44 392 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=52780 $D=0
M2093 203 44 393 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=57410 $D=0
M2094 204 44 394 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=62040 $D=0
M2095 205 44 395 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=66670 $D=0
M2096 396 45 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=52780 $D=0
M2097 397 45 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=57410 $D=0
M2098 398 45 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=62040 $D=0
M2099 399 45 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=66670 $D=0
M2100 400 392 280 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=52780 $D=0
M2101 401 393 281 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=57410 $D=0
M2102 402 394 282 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=62040 $D=0
M2103 403 395 283 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=66670 $D=0
M2104 202 400 1254 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=52780 $D=0
M2105 203 401 1255 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=57410 $D=0
M2106 204 402 1256 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=62040 $D=0
M2107 205 403 1257 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=66670 $D=0
M2108 404 1254 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=52780 $D=0
M2109 405 1255 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=57410 $D=0
M2110 406 1256 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=62040 $D=0
M2111 407 1257 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=66670 $D=0
M2112 400 44 404 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=52780 $D=0
M2113 401 44 405 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=57410 $D=0
M2114 402 44 406 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=62040 $D=0
M2115 403 44 407 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=66670 $D=0
M2116 404 396 300 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=52780 $D=0
M2117 405 397 301 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=57410 $D=0
M2118 406 398 302 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=62040 $D=0
M2119 407 399 303 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=66670 $D=0
M2120 308 408 404 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=52780 $D=0
M2121 309 409 405 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=57410 $D=0
M2122 310 410 406 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=62040 $D=0
M2123 311 411 407 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=66670 $D=0
M2124 408 46 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=52780 $D=0
M2125 409 46 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=57410 $D=0
M2126 410 46 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=62040 $D=0
M2127 411 46 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=66670 $D=0
M2128 202 47 412 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=52780 $D=0
M2129 203 47 413 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=57410 $D=0
M2130 204 47 414 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=62040 $D=0
M2131 205 47 415 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=66670 $D=0
M2132 416 48 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=52780 $D=0
M2133 417 48 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=57410 $D=0
M2134 418 48 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=62040 $D=0
M2135 419 48 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=66670 $D=0
M2136 420 412 280 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=52780 $D=0
M2137 421 413 281 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=57410 $D=0
M2138 422 414 282 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=62040 $D=0
M2139 423 415 283 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=66670 $D=0
M2140 202 420 1258 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=52780 $D=0
M2141 203 421 1259 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=57410 $D=0
M2142 204 422 1260 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=62040 $D=0
M2143 205 423 1261 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=66670 $D=0
M2144 424 1258 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=52780 $D=0
M2145 425 1259 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=57410 $D=0
M2146 426 1260 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=62040 $D=0
M2147 427 1261 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=66670 $D=0
M2148 420 47 424 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=52780 $D=0
M2149 421 47 425 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=57410 $D=0
M2150 422 47 426 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=62040 $D=0
M2151 423 47 427 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=66670 $D=0
M2152 424 416 300 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=52780 $D=0
M2153 425 417 301 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=57410 $D=0
M2154 426 418 302 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=62040 $D=0
M2155 427 419 303 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=66670 $D=0
M2156 308 428 424 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=52780 $D=0
M2157 309 429 425 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=57410 $D=0
M2158 310 430 426 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=62040 $D=0
M2159 311 431 427 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=66670 $D=0
M2160 428 49 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=52780 $D=0
M2161 429 49 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=57410 $D=0
M2162 430 49 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=62040 $D=0
M2163 431 49 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=66670 $D=0
M2164 202 50 432 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=52780 $D=0
M2165 203 50 433 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=57410 $D=0
M2166 204 50 434 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=62040 $D=0
M2167 205 50 435 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=66670 $D=0
M2168 436 51 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=52780 $D=0
M2169 437 51 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=57410 $D=0
M2170 438 51 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=62040 $D=0
M2171 439 51 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=66670 $D=0
M2172 440 432 280 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=52780 $D=0
M2173 441 433 281 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=57410 $D=0
M2174 442 434 282 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=62040 $D=0
M2175 443 435 283 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=66670 $D=0
M2176 202 440 1262 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=52780 $D=0
M2177 203 441 1263 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=57410 $D=0
M2178 204 442 1264 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=62040 $D=0
M2179 205 443 1265 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=66670 $D=0
M2180 444 1262 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=52780 $D=0
M2181 445 1263 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=57410 $D=0
M2182 446 1264 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=62040 $D=0
M2183 447 1265 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=66670 $D=0
M2184 440 50 444 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=52780 $D=0
M2185 441 50 445 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=57410 $D=0
M2186 442 50 446 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=62040 $D=0
M2187 443 50 447 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=66670 $D=0
M2188 444 436 300 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=52780 $D=0
M2189 445 437 301 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=57410 $D=0
M2190 446 438 302 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=62040 $D=0
M2191 447 439 303 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=66670 $D=0
M2192 308 448 444 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=52780 $D=0
M2193 309 449 445 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=57410 $D=0
M2194 310 450 446 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=62040 $D=0
M2195 311 451 447 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=66670 $D=0
M2196 448 52 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=52780 $D=0
M2197 449 52 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=57410 $D=0
M2198 450 52 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=62040 $D=0
M2199 451 52 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=66670 $D=0
M2200 202 53 452 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=52780 $D=0
M2201 203 53 453 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=57410 $D=0
M2202 204 53 454 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=62040 $D=0
M2203 205 53 455 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=66670 $D=0
M2204 456 54 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=52780 $D=0
M2205 457 54 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=57410 $D=0
M2206 458 54 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=62040 $D=0
M2207 459 54 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=66670 $D=0
M2208 460 452 280 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=52780 $D=0
M2209 461 453 281 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=57410 $D=0
M2210 462 454 282 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=62040 $D=0
M2211 463 455 283 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=66670 $D=0
M2212 202 460 1266 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=52780 $D=0
M2213 203 461 1267 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=57410 $D=0
M2214 204 462 1268 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=62040 $D=0
M2215 205 463 1269 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=66670 $D=0
M2216 464 1266 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=52780 $D=0
M2217 465 1267 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=57410 $D=0
M2218 466 1268 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=62040 $D=0
M2219 467 1269 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=66670 $D=0
M2220 460 53 464 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=52780 $D=0
M2221 461 53 465 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=57410 $D=0
M2222 462 53 466 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=62040 $D=0
M2223 463 53 467 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=66670 $D=0
M2224 464 456 300 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=52780 $D=0
M2225 465 457 301 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=57410 $D=0
M2226 466 458 302 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=62040 $D=0
M2227 467 459 303 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=66670 $D=0
M2228 308 468 464 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=52780 $D=0
M2229 309 469 465 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=57410 $D=0
M2230 310 470 466 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=62040 $D=0
M2231 311 471 467 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=66670 $D=0
M2232 468 55 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=52780 $D=0
M2233 469 55 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=57410 $D=0
M2234 470 55 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=62040 $D=0
M2235 471 55 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=66670 $D=0
M2236 202 56 472 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=52780 $D=0
M2237 203 56 473 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=57410 $D=0
M2238 204 56 474 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=62040 $D=0
M2239 205 56 475 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=66670 $D=0
M2240 476 57 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=52780 $D=0
M2241 477 57 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=57410 $D=0
M2242 478 57 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=62040 $D=0
M2243 479 57 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=66670 $D=0
M2244 480 472 280 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=52780 $D=0
M2245 481 473 281 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=57410 $D=0
M2246 482 474 282 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=62040 $D=0
M2247 483 475 283 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=66670 $D=0
M2248 202 480 1270 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=52780 $D=0
M2249 203 481 1271 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=57410 $D=0
M2250 204 482 1272 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=62040 $D=0
M2251 205 483 1273 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=66670 $D=0
M2252 484 1270 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=52780 $D=0
M2253 485 1271 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=57410 $D=0
M2254 486 1272 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=62040 $D=0
M2255 487 1273 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=66670 $D=0
M2256 480 56 484 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=52780 $D=0
M2257 481 56 485 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=57410 $D=0
M2258 482 56 486 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=62040 $D=0
M2259 483 56 487 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=66670 $D=0
M2260 484 476 300 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=52780 $D=0
M2261 485 477 301 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=57410 $D=0
M2262 486 478 302 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=62040 $D=0
M2263 487 479 303 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=66670 $D=0
M2264 308 488 484 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=52780 $D=0
M2265 309 489 485 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=57410 $D=0
M2266 310 490 486 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=62040 $D=0
M2267 311 491 487 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=66670 $D=0
M2268 488 58 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=52780 $D=0
M2269 489 58 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=57410 $D=0
M2270 490 58 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=62040 $D=0
M2271 491 58 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=66670 $D=0
M2272 202 59 492 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=52780 $D=0
M2273 203 59 493 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=57410 $D=0
M2274 204 59 494 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=62040 $D=0
M2275 205 59 495 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=66670 $D=0
M2276 496 60 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=52780 $D=0
M2277 497 60 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=57410 $D=0
M2278 498 60 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=62040 $D=0
M2279 499 60 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=66670 $D=0
M2280 500 492 280 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=52780 $D=0
M2281 501 493 281 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=57410 $D=0
M2282 502 494 282 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=62040 $D=0
M2283 503 495 283 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=66670 $D=0
M2284 202 500 1274 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=52780 $D=0
M2285 203 501 1275 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=57410 $D=0
M2286 204 502 1276 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=62040 $D=0
M2287 205 503 1277 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=66670 $D=0
M2288 504 1274 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=52780 $D=0
M2289 505 1275 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=57410 $D=0
M2290 506 1276 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=62040 $D=0
M2291 507 1277 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=66670 $D=0
M2292 500 59 504 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=52780 $D=0
M2293 501 59 505 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=57410 $D=0
M2294 502 59 506 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=62040 $D=0
M2295 503 59 507 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=66670 $D=0
M2296 504 496 300 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=52780 $D=0
M2297 505 497 301 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=57410 $D=0
M2298 506 498 302 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=62040 $D=0
M2299 507 499 303 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=66670 $D=0
M2300 308 508 504 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=52780 $D=0
M2301 309 509 505 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=57410 $D=0
M2302 310 510 506 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=62040 $D=0
M2303 311 511 507 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=66670 $D=0
M2304 508 61 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=52780 $D=0
M2305 509 61 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=57410 $D=0
M2306 510 61 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=62040 $D=0
M2307 511 61 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=66670 $D=0
M2308 202 62 512 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=52780 $D=0
M2309 203 62 513 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=57410 $D=0
M2310 204 62 514 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=62040 $D=0
M2311 205 62 515 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=66670 $D=0
M2312 516 63 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=52780 $D=0
M2313 517 63 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=57410 $D=0
M2314 518 63 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=62040 $D=0
M2315 519 63 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=66670 $D=0
M2316 520 512 280 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=52780 $D=0
M2317 521 513 281 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=57410 $D=0
M2318 522 514 282 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=62040 $D=0
M2319 523 515 283 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=66670 $D=0
M2320 202 520 1278 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=52780 $D=0
M2321 203 521 1279 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=57410 $D=0
M2322 204 522 1280 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=62040 $D=0
M2323 205 523 1281 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=66670 $D=0
M2324 524 1278 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=52780 $D=0
M2325 525 1279 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=57410 $D=0
M2326 526 1280 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=62040 $D=0
M2327 527 1281 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=66670 $D=0
M2328 520 62 524 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=52780 $D=0
M2329 521 62 525 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=57410 $D=0
M2330 522 62 526 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=62040 $D=0
M2331 523 62 527 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=66670 $D=0
M2332 524 516 300 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=52780 $D=0
M2333 525 517 301 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=57410 $D=0
M2334 526 518 302 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=62040 $D=0
M2335 527 519 303 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=66670 $D=0
M2336 308 528 524 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=52780 $D=0
M2337 309 529 525 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=57410 $D=0
M2338 310 530 526 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=62040 $D=0
M2339 311 531 527 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=66670 $D=0
M2340 528 64 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=52780 $D=0
M2341 529 64 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=57410 $D=0
M2342 530 64 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=62040 $D=0
M2343 531 64 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=66670 $D=0
M2344 202 65 532 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=52780 $D=0
M2345 203 65 533 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=57410 $D=0
M2346 204 65 534 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=62040 $D=0
M2347 205 65 535 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=66670 $D=0
M2348 536 66 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=52780 $D=0
M2349 537 66 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=57410 $D=0
M2350 538 66 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=62040 $D=0
M2351 539 66 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=66670 $D=0
M2352 540 532 280 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=52780 $D=0
M2353 541 533 281 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=57410 $D=0
M2354 542 534 282 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=62040 $D=0
M2355 543 535 283 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=66670 $D=0
M2356 202 540 1282 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=52780 $D=0
M2357 203 541 1283 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=57410 $D=0
M2358 204 542 1284 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=62040 $D=0
M2359 205 543 1285 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=66670 $D=0
M2360 544 1282 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=52780 $D=0
M2361 545 1283 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=57410 $D=0
M2362 546 1284 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=62040 $D=0
M2363 547 1285 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=66670 $D=0
M2364 540 65 544 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=52780 $D=0
M2365 541 65 545 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=57410 $D=0
M2366 542 65 546 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=62040 $D=0
M2367 543 65 547 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=66670 $D=0
M2368 544 536 300 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=52780 $D=0
M2369 545 537 301 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=57410 $D=0
M2370 546 538 302 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=62040 $D=0
M2371 547 539 303 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=66670 $D=0
M2372 308 548 544 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=52780 $D=0
M2373 309 549 545 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=57410 $D=0
M2374 310 550 546 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=62040 $D=0
M2375 311 551 547 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=66670 $D=0
M2376 548 67 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=52780 $D=0
M2377 549 67 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=57410 $D=0
M2378 550 67 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=62040 $D=0
M2379 551 67 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=66670 $D=0
M2380 202 68 552 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=52780 $D=0
M2381 203 68 553 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=57410 $D=0
M2382 204 68 554 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=62040 $D=0
M2383 205 68 555 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=66670 $D=0
M2384 556 69 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=52780 $D=0
M2385 557 69 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=57410 $D=0
M2386 558 69 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=62040 $D=0
M2387 559 69 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=66670 $D=0
M2388 560 552 280 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=52780 $D=0
M2389 561 553 281 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=57410 $D=0
M2390 562 554 282 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=62040 $D=0
M2391 563 555 283 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=66670 $D=0
M2392 202 560 1286 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=52780 $D=0
M2393 203 561 1287 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=57410 $D=0
M2394 204 562 1288 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=62040 $D=0
M2395 205 563 1289 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=66670 $D=0
M2396 564 1286 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=52780 $D=0
M2397 565 1287 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=57410 $D=0
M2398 566 1288 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=62040 $D=0
M2399 567 1289 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=66670 $D=0
M2400 560 68 564 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=52780 $D=0
M2401 561 68 565 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=57410 $D=0
M2402 562 68 566 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=62040 $D=0
M2403 563 68 567 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=66670 $D=0
M2404 564 556 300 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=52780 $D=0
M2405 565 557 301 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=57410 $D=0
M2406 566 558 302 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=62040 $D=0
M2407 567 559 303 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=66670 $D=0
M2408 308 568 564 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=52780 $D=0
M2409 309 569 565 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=57410 $D=0
M2410 310 570 566 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=62040 $D=0
M2411 311 571 567 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=66670 $D=0
M2412 568 70 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=52780 $D=0
M2413 569 70 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=57410 $D=0
M2414 570 70 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=62040 $D=0
M2415 571 70 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=66670 $D=0
M2416 202 71 572 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=52780 $D=0
M2417 203 71 573 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=57410 $D=0
M2418 204 71 574 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=62040 $D=0
M2419 205 71 575 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=66670 $D=0
M2420 576 72 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=52780 $D=0
M2421 577 72 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=57410 $D=0
M2422 578 72 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=62040 $D=0
M2423 579 72 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=66670 $D=0
M2424 580 572 280 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=52780 $D=0
M2425 581 573 281 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=57410 $D=0
M2426 582 574 282 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=62040 $D=0
M2427 583 575 283 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=66670 $D=0
M2428 202 580 1290 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=52780 $D=0
M2429 203 581 1291 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=57410 $D=0
M2430 204 582 1292 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=62040 $D=0
M2431 205 583 1293 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=66670 $D=0
M2432 584 1290 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=52780 $D=0
M2433 585 1291 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=57410 $D=0
M2434 586 1292 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=62040 $D=0
M2435 587 1293 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=66670 $D=0
M2436 580 71 584 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=52780 $D=0
M2437 581 71 585 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=57410 $D=0
M2438 582 71 586 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=62040 $D=0
M2439 583 71 587 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=66670 $D=0
M2440 584 576 300 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=52780 $D=0
M2441 585 577 301 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=57410 $D=0
M2442 586 578 302 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=62040 $D=0
M2443 587 579 303 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=66670 $D=0
M2444 308 588 584 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=52780 $D=0
M2445 309 589 585 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=57410 $D=0
M2446 310 590 586 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=62040 $D=0
M2447 311 591 587 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=66670 $D=0
M2448 588 73 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=52780 $D=0
M2449 589 73 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=57410 $D=0
M2450 590 73 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=62040 $D=0
M2451 591 73 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=66670 $D=0
M2452 202 74 592 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=52780 $D=0
M2453 203 74 593 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=57410 $D=0
M2454 204 74 594 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=62040 $D=0
M2455 205 74 595 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=66670 $D=0
M2456 596 75 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=52780 $D=0
M2457 597 75 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=57410 $D=0
M2458 598 75 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=62040 $D=0
M2459 599 75 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=66670 $D=0
M2460 600 592 280 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=52780 $D=0
M2461 601 593 281 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=57410 $D=0
M2462 602 594 282 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=62040 $D=0
M2463 603 595 283 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=66670 $D=0
M2464 202 600 1294 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=52780 $D=0
M2465 203 601 1295 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=57410 $D=0
M2466 204 602 1296 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=62040 $D=0
M2467 205 603 1297 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=66670 $D=0
M2468 604 1294 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=52780 $D=0
M2469 605 1295 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=57410 $D=0
M2470 606 1296 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=62040 $D=0
M2471 607 1297 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=66670 $D=0
M2472 600 74 604 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=52780 $D=0
M2473 601 74 605 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=57410 $D=0
M2474 602 74 606 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=62040 $D=0
M2475 603 74 607 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=66670 $D=0
M2476 604 596 300 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=52780 $D=0
M2477 605 597 301 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=57410 $D=0
M2478 606 598 302 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=62040 $D=0
M2479 607 599 303 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=66670 $D=0
M2480 308 608 604 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=52780 $D=0
M2481 309 609 605 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=57410 $D=0
M2482 310 610 606 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=62040 $D=0
M2483 311 611 607 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=66670 $D=0
M2484 608 76 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=52780 $D=0
M2485 609 76 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=57410 $D=0
M2486 610 76 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=62040 $D=0
M2487 611 76 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=66670 $D=0
M2488 202 77 612 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=52780 $D=0
M2489 203 77 613 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=57410 $D=0
M2490 204 77 614 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=62040 $D=0
M2491 205 77 615 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=66670 $D=0
M2492 616 78 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=52780 $D=0
M2493 617 78 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=57410 $D=0
M2494 618 78 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=62040 $D=0
M2495 619 78 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=66670 $D=0
M2496 620 612 280 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=52780 $D=0
M2497 621 613 281 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=57410 $D=0
M2498 622 614 282 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=62040 $D=0
M2499 623 615 283 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=66670 $D=0
M2500 202 620 1298 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=52780 $D=0
M2501 203 621 1299 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=57410 $D=0
M2502 204 622 1300 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=62040 $D=0
M2503 205 623 1301 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=66670 $D=0
M2504 624 1298 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=52780 $D=0
M2505 625 1299 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=57410 $D=0
M2506 626 1300 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=62040 $D=0
M2507 627 1301 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=66670 $D=0
M2508 620 77 624 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=52780 $D=0
M2509 621 77 625 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=57410 $D=0
M2510 622 77 626 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=62040 $D=0
M2511 623 77 627 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=66670 $D=0
M2512 624 616 300 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=52780 $D=0
M2513 625 617 301 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=57410 $D=0
M2514 626 618 302 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=62040 $D=0
M2515 627 619 303 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=66670 $D=0
M2516 308 628 624 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=52780 $D=0
M2517 309 629 625 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=57410 $D=0
M2518 310 630 626 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=62040 $D=0
M2519 311 631 627 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=66670 $D=0
M2520 628 79 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=52780 $D=0
M2521 629 79 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=57410 $D=0
M2522 630 79 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=62040 $D=0
M2523 631 79 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=66670 $D=0
M2524 202 80 632 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=52780 $D=0
M2525 203 80 633 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=57410 $D=0
M2526 204 80 634 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=62040 $D=0
M2527 205 80 635 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=66670 $D=0
M2528 636 81 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=52780 $D=0
M2529 637 81 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=57410 $D=0
M2530 638 81 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=62040 $D=0
M2531 639 81 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=66670 $D=0
M2532 640 632 280 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=52780 $D=0
M2533 641 633 281 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=57410 $D=0
M2534 642 634 282 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=62040 $D=0
M2535 643 635 283 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=66670 $D=0
M2536 202 640 1302 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=52780 $D=0
M2537 203 641 1303 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=57410 $D=0
M2538 204 642 1304 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=62040 $D=0
M2539 205 643 1305 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=66670 $D=0
M2540 644 1302 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=52780 $D=0
M2541 645 1303 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=57410 $D=0
M2542 646 1304 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=62040 $D=0
M2543 647 1305 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=66670 $D=0
M2544 640 80 644 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=52780 $D=0
M2545 641 80 645 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=57410 $D=0
M2546 642 80 646 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=62040 $D=0
M2547 643 80 647 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=66670 $D=0
M2548 644 636 300 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=52780 $D=0
M2549 645 637 301 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=57410 $D=0
M2550 646 638 302 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=62040 $D=0
M2551 647 639 303 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=66670 $D=0
M2552 308 648 644 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=52780 $D=0
M2553 309 649 645 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=57410 $D=0
M2554 310 650 646 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=62040 $D=0
M2555 311 651 647 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=66670 $D=0
M2556 648 82 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=52780 $D=0
M2557 649 82 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=57410 $D=0
M2558 650 82 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=62040 $D=0
M2559 651 82 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=66670 $D=0
M2560 202 83 652 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=52780 $D=0
M2561 203 83 653 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=57410 $D=0
M2562 204 83 654 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=62040 $D=0
M2563 205 83 655 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=66670 $D=0
M2564 656 84 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=52780 $D=0
M2565 657 84 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=57410 $D=0
M2566 658 84 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=62040 $D=0
M2567 659 84 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=66670 $D=0
M2568 660 652 280 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=52780 $D=0
M2569 661 653 281 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=57410 $D=0
M2570 662 654 282 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=62040 $D=0
M2571 663 655 283 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=66670 $D=0
M2572 202 660 1306 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=52780 $D=0
M2573 203 661 1307 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=57410 $D=0
M2574 204 662 1308 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=62040 $D=0
M2575 205 663 1309 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=66670 $D=0
M2576 664 1306 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=52780 $D=0
M2577 665 1307 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=57410 $D=0
M2578 666 1308 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=62040 $D=0
M2579 667 1309 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=66670 $D=0
M2580 660 83 664 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=52780 $D=0
M2581 661 83 665 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=57410 $D=0
M2582 662 83 666 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=62040 $D=0
M2583 663 83 667 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=66670 $D=0
M2584 664 656 300 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=52780 $D=0
M2585 665 657 301 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=57410 $D=0
M2586 666 658 302 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=62040 $D=0
M2587 667 659 303 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=66670 $D=0
M2588 308 668 664 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=52780 $D=0
M2589 309 669 665 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=57410 $D=0
M2590 310 670 666 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=62040 $D=0
M2591 311 671 667 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=66670 $D=0
M2592 668 85 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=52780 $D=0
M2593 669 85 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=57410 $D=0
M2594 670 85 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=62040 $D=0
M2595 671 85 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=66670 $D=0
M2596 202 86 672 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=52780 $D=0
M2597 203 86 673 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=57410 $D=0
M2598 204 86 674 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=62040 $D=0
M2599 205 86 675 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=66670 $D=0
M2600 676 87 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=52780 $D=0
M2601 677 87 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=57410 $D=0
M2602 678 87 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=62040 $D=0
M2603 679 87 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=66670 $D=0
M2604 680 672 280 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=52780 $D=0
M2605 681 673 281 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=57410 $D=0
M2606 682 674 282 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=62040 $D=0
M2607 683 675 283 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=66670 $D=0
M2608 202 680 1310 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=52780 $D=0
M2609 203 681 1311 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=57410 $D=0
M2610 204 682 1312 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=62040 $D=0
M2611 205 683 1313 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=66670 $D=0
M2612 684 1310 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=52780 $D=0
M2613 685 1311 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=57410 $D=0
M2614 686 1312 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=62040 $D=0
M2615 687 1313 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=66670 $D=0
M2616 680 86 684 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=52780 $D=0
M2617 681 86 685 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=57410 $D=0
M2618 682 86 686 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=62040 $D=0
M2619 683 86 687 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=66670 $D=0
M2620 684 676 300 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=52780 $D=0
M2621 685 677 301 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=57410 $D=0
M2622 686 678 302 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=62040 $D=0
M2623 687 679 303 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=66670 $D=0
M2624 308 688 684 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=52780 $D=0
M2625 309 689 685 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=57410 $D=0
M2626 310 690 686 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=62040 $D=0
M2627 311 691 687 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=66670 $D=0
M2628 688 88 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=52780 $D=0
M2629 689 88 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=57410 $D=0
M2630 690 88 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=62040 $D=0
M2631 691 88 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=66670 $D=0
M2632 202 89 692 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=52780 $D=0
M2633 203 89 693 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=57410 $D=0
M2634 204 89 694 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=62040 $D=0
M2635 205 89 695 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=66670 $D=0
M2636 696 90 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=52780 $D=0
M2637 697 90 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=57410 $D=0
M2638 698 90 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=62040 $D=0
M2639 699 90 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=66670 $D=0
M2640 700 692 280 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=52780 $D=0
M2641 701 693 281 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=57410 $D=0
M2642 702 694 282 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=62040 $D=0
M2643 703 695 283 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=66670 $D=0
M2644 202 700 1314 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=52780 $D=0
M2645 203 701 1315 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=57410 $D=0
M2646 204 702 1316 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=62040 $D=0
M2647 205 703 1317 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=66670 $D=0
M2648 704 1314 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=52780 $D=0
M2649 705 1315 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=57410 $D=0
M2650 706 1316 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=62040 $D=0
M2651 707 1317 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=66670 $D=0
M2652 700 89 704 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=52780 $D=0
M2653 701 89 705 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=57410 $D=0
M2654 702 89 706 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=62040 $D=0
M2655 703 89 707 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=66670 $D=0
M2656 704 696 300 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=52780 $D=0
M2657 705 697 301 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=57410 $D=0
M2658 706 698 302 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=62040 $D=0
M2659 707 699 303 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=66670 $D=0
M2660 308 708 704 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=52780 $D=0
M2661 309 709 705 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=57410 $D=0
M2662 310 710 706 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=62040 $D=0
M2663 311 711 707 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=66670 $D=0
M2664 708 91 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=52780 $D=0
M2665 709 91 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=57410 $D=0
M2666 710 91 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=62040 $D=0
M2667 711 91 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=66670 $D=0
M2668 202 92 712 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=52780 $D=0
M2669 203 92 713 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=57410 $D=0
M2670 204 92 714 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=62040 $D=0
M2671 205 92 715 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=66670 $D=0
M2672 716 93 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=52780 $D=0
M2673 717 93 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=57410 $D=0
M2674 718 93 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=62040 $D=0
M2675 719 93 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=66670 $D=0
M2676 720 712 280 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=52780 $D=0
M2677 721 713 281 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=57410 $D=0
M2678 722 714 282 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=62040 $D=0
M2679 723 715 283 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=66670 $D=0
M2680 202 720 1318 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=52780 $D=0
M2681 203 721 1319 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=57410 $D=0
M2682 204 722 1320 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=62040 $D=0
M2683 205 723 1321 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=66670 $D=0
M2684 724 1318 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=52780 $D=0
M2685 725 1319 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=57410 $D=0
M2686 726 1320 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=62040 $D=0
M2687 727 1321 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=66670 $D=0
M2688 720 92 724 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=52780 $D=0
M2689 721 92 725 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=57410 $D=0
M2690 722 92 726 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=62040 $D=0
M2691 723 92 727 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=66670 $D=0
M2692 724 716 300 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=52780 $D=0
M2693 725 717 301 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=57410 $D=0
M2694 726 718 302 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=62040 $D=0
M2695 727 719 303 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=66670 $D=0
M2696 308 728 724 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=52780 $D=0
M2697 309 729 725 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=57410 $D=0
M2698 310 730 726 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=62040 $D=0
M2699 311 731 727 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=66670 $D=0
M2700 728 94 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=52780 $D=0
M2701 729 94 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=57410 $D=0
M2702 730 94 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=62040 $D=0
M2703 731 94 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=66670 $D=0
M2704 202 95 732 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=52780 $D=0
M2705 203 95 733 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=57410 $D=0
M2706 204 95 734 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=62040 $D=0
M2707 205 95 735 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=66670 $D=0
M2708 736 96 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=52780 $D=0
M2709 737 96 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=57410 $D=0
M2710 738 96 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=62040 $D=0
M2711 739 96 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=66670 $D=0
M2712 740 732 280 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=52780 $D=0
M2713 741 733 281 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=57410 $D=0
M2714 742 734 282 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=62040 $D=0
M2715 743 735 283 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=66670 $D=0
M2716 202 740 1322 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=52780 $D=0
M2717 203 741 1323 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=57410 $D=0
M2718 204 742 1324 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=62040 $D=0
M2719 205 743 1325 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=66670 $D=0
M2720 744 1322 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=52780 $D=0
M2721 745 1323 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=57410 $D=0
M2722 746 1324 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=62040 $D=0
M2723 747 1325 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=66670 $D=0
M2724 740 95 744 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=52780 $D=0
M2725 741 95 745 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=57410 $D=0
M2726 742 95 746 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=62040 $D=0
M2727 743 95 747 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=66670 $D=0
M2728 744 736 300 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=52780 $D=0
M2729 745 737 301 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=57410 $D=0
M2730 746 738 302 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=62040 $D=0
M2731 747 739 303 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=66670 $D=0
M2732 308 748 744 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=52780 $D=0
M2733 309 749 745 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=57410 $D=0
M2734 310 750 746 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=62040 $D=0
M2735 311 751 747 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=66670 $D=0
M2736 748 97 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=52780 $D=0
M2737 749 97 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=57410 $D=0
M2738 750 97 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=62040 $D=0
M2739 751 97 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=66670 $D=0
M2740 202 98 752 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=52780 $D=0
M2741 203 98 753 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=57410 $D=0
M2742 204 98 754 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=62040 $D=0
M2743 205 98 755 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=66670 $D=0
M2744 756 99 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=52780 $D=0
M2745 757 99 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=57410 $D=0
M2746 758 99 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=62040 $D=0
M2747 759 99 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=66670 $D=0
M2748 760 752 280 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=52780 $D=0
M2749 761 753 281 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=57410 $D=0
M2750 762 754 282 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=62040 $D=0
M2751 763 755 283 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=66670 $D=0
M2752 202 760 1326 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=52780 $D=0
M2753 203 761 1327 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=57410 $D=0
M2754 204 762 1328 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=62040 $D=0
M2755 205 763 1329 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=66670 $D=0
M2756 764 1326 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=52780 $D=0
M2757 765 1327 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=57410 $D=0
M2758 766 1328 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=62040 $D=0
M2759 767 1329 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=66670 $D=0
M2760 760 98 764 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=52780 $D=0
M2761 761 98 765 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=57410 $D=0
M2762 762 98 766 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=62040 $D=0
M2763 763 98 767 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=66670 $D=0
M2764 764 756 300 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=52780 $D=0
M2765 765 757 301 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=57410 $D=0
M2766 766 758 302 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=62040 $D=0
M2767 767 759 303 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=66670 $D=0
M2768 308 768 764 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=52780 $D=0
M2769 309 769 765 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=57410 $D=0
M2770 310 770 766 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=62040 $D=0
M2771 311 771 767 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=66670 $D=0
M2772 768 100 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=52780 $D=0
M2773 769 100 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=57410 $D=0
M2774 770 100 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=62040 $D=0
M2775 771 100 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=66670 $D=0
M2776 202 101 772 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=52780 $D=0
M2777 203 101 773 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=57410 $D=0
M2778 204 101 774 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=62040 $D=0
M2779 205 101 775 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=66670 $D=0
M2780 776 102 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=52780 $D=0
M2781 777 102 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=57410 $D=0
M2782 778 102 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=62040 $D=0
M2783 779 102 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=66670 $D=0
M2784 780 772 280 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=52780 $D=0
M2785 781 773 281 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=57410 $D=0
M2786 782 774 282 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=62040 $D=0
M2787 783 775 283 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=66670 $D=0
M2788 202 780 1330 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=52780 $D=0
M2789 203 781 1331 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=57410 $D=0
M2790 204 782 1332 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=62040 $D=0
M2791 205 783 1333 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=66670 $D=0
M2792 784 1330 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=52780 $D=0
M2793 785 1331 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=57410 $D=0
M2794 786 1332 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=62040 $D=0
M2795 787 1333 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=66670 $D=0
M2796 780 101 784 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=52780 $D=0
M2797 781 101 785 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=57410 $D=0
M2798 782 101 786 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=62040 $D=0
M2799 783 101 787 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=66670 $D=0
M2800 784 776 300 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=52780 $D=0
M2801 785 777 301 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=57410 $D=0
M2802 786 778 302 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=62040 $D=0
M2803 787 779 303 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=66670 $D=0
M2804 308 788 784 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=52780 $D=0
M2805 309 789 785 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=57410 $D=0
M2806 310 790 786 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=62040 $D=0
M2807 311 791 787 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=66670 $D=0
M2808 788 103 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=52780 $D=0
M2809 789 103 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=57410 $D=0
M2810 790 103 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=62040 $D=0
M2811 791 103 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=66670 $D=0
M2812 202 104 792 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=52780 $D=0
M2813 203 104 793 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=57410 $D=0
M2814 204 104 794 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=62040 $D=0
M2815 205 104 795 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=66670 $D=0
M2816 796 105 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=52780 $D=0
M2817 797 105 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=57410 $D=0
M2818 798 105 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=62040 $D=0
M2819 799 105 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=66670 $D=0
M2820 800 792 280 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=52780 $D=0
M2821 801 793 281 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=57410 $D=0
M2822 802 794 282 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=62040 $D=0
M2823 803 795 283 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=66670 $D=0
M2824 202 800 1334 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=52780 $D=0
M2825 203 801 1335 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=57410 $D=0
M2826 204 802 1336 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=62040 $D=0
M2827 205 803 1337 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=66670 $D=0
M2828 804 1334 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=52780 $D=0
M2829 805 1335 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=57410 $D=0
M2830 806 1336 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=62040 $D=0
M2831 807 1337 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=66670 $D=0
M2832 800 104 804 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=52780 $D=0
M2833 801 104 805 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=57410 $D=0
M2834 802 104 806 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=62040 $D=0
M2835 803 104 807 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=66670 $D=0
M2836 804 796 300 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=52780 $D=0
M2837 805 797 301 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=57410 $D=0
M2838 806 798 302 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=62040 $D=0
M2839 807 799 303 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=66670 $D=0
M2840 308 808 804 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=52780 $D=0
M2841 309 809 805 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=57410 $D=0
M2842 310 810 806 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=62040 $D=0
M2843 311 811 807 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=66670 $D=0
M2844 808 106 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=52780 $D=0
M2845 809 106 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=57410 $D=0
M2846 810 106 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=62040 $D=0
M2847 811 106 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=66670 $D=0
M2848 202 107 812 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=52780 $D=0
M2849 203 107 813 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=57410 $D=0
M2850 204 107 814 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=62040 $D=0
M2851 205 107 815 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=66670 $D=0
M2852 816 108 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=52780 $D=0
M2853 817 108 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=57410 $D=0
M2854 818 108 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=62040 $D=0
M2855 819 108 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=66670 $D=0
M2856 820 812 280 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=52780 $D=0
M2857 821 813 281 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=57410 $D=0
M2858 822 814 282 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=62040 $D=0
M2859 823 815 283 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=66670 $D=0
M2860 202 820 1338 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=52780 $D=0
M2861 203 821 1339 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=57410 $D=0
M2862 204 822 1340 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=62040 $D=0
M2863 205 823 1341 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=66670 $D=0
M2864 824 1338 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=52780 $D=0
M2865 825 1339 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=57410 $D=0
M2866 826 1340 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=62040 $D=0
M2867 827 1341 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=66670 $D=0
M2868 820 107 824 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=52780 $D=0
M2869 821 107 825 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=57410 $D=0
M2870 822 107 826 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=62040 $D=0
M2871 823 107 827 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=66670 $D=0
M2872 824 816 300 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=52780 $D=0
M2873 825 817 301 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=57410 $D=0
M2874 826 818 302 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=62040 $D=0
M2875 827 819 303 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=66670 $D=0
M2876 308 828 824 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=52780 $D=0
M2877 309 829 825 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=57410 $D=0
M2878 310 830 826 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=62040 $D=0
M2879 311 831 827 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=66670 $D=0
M2880 828 109 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=52780 $D=0
M2881 829 109 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=57410 $D=0
M2882 830 109 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=62040 $D=0
M2883 831 109 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=66670 $D=0
M2884 202 110 832 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=52780 $D=0
M2885 203 110 833 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=57410 $D=0
M2886 204 110 834 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=62040 $D=0
M2887 205 110 835 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=66670 $D=0
M2888 836 111 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=52780 $D=0
M2889 837 111 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=57410 $D=0
M2890 838 111 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=62040 $D=0
M2891 839 111 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=66670 $D=0
M2892 840 832 280 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=52780 $D=0
M2893 841 833 281 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=57410 $D=0
M2894 842 834 282 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=62040 $D=0
M2895 843 835 283 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=66670 $D=0
M2896 202 840 1342 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=52780 $D=0
M2897 203 841 1343 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=57410 $D=0
M2898 204 842 1344 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=62040 $D=0
M2899 205 843 1345 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=66670 $D=0
M2900 844 1342 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=52780 $D=0
M2901 845 1343 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=57410 $D=0
M2902 846 1344 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=62040 $D=0
M2903 847 1345 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=66670 $D=0
M2904 840 110 844 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=52780 $D=0
M2905 841 110 845 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=57410 $D=0
M2906 842 110 846 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=62040 $D=0
M2907 843 110 847 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=66670 $D=0
M2908 844 836 300 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=52780 $D=0
M2909 845 837 301 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=57410 $D=0
M2910 846 838 302 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=62040 $D=0
M2911 847 839 303 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=66670 $D=0
M2912 308 848 844 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=52780 $D=0
M2913 309 849 845 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=57410 $D=0
M2914 310 850 846 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=62040 $D=0
M2915 311 851 847 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=66670 $D=0
M2916 848 112 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=52780 $D=0
M2917 849 112 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=57410 $D=0
M2918 850 112 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=62040 $D=0
M2919 851 112 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=66670 $D=0
M2920 202 113 852 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=52780 $D=0
M2921 203 113 853 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=57410 $D=0
M2922 204 113 854 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=62040 $D=0
M2923 205 113 855 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=66670 $D=0
M2924 856 114 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=52780 $D=0
M2925 857 114 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=57410 $D=0
M2926 858 114 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=62040 $D=0
M2927 859 114 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=66670 $D=0
M2928 860 852 280 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=52780 $D=0
M2929 861 853 281 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=57410 $D=0
M2930 862 854 282 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=62040 $D=0
M2931 863 855 283 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=66670 $D=0
M2932 202 860 1346 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=52780 $D=0
M2933 203 861 1347 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=57410 $D=0
M2934 204 862 1348 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=62040 $D=0
M2935 205 863 1349 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=66670 $D=0
M2936 864 1346 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=52780 $D=0
M2937 865 1347 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=57410 $D=0
M2938 866 1348 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=62040 $D=0
M2939 867 1349 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=66670 $D=0
M2940 860 113 864 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=52780 $D=0
M2941 861 113 865 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=57410 $D=0
M2942 862 113 866 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=62040 $D=0
M2943 863 113 867 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=66670 $D=0
M2944 864 856 300 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=52780 $D=0
M2945 865 857 301 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=57410 $D=0
M2946 866 858 302 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=62040 $D=0
M2947 867 859 303 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=66670 $D=0
M2948 308 868 864 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=52780 $D=0
M2949 309 869 865 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=57410 $D=0
M2950 310 870 866 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=62040 $D=0
M2951 311 871 867 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=66670 $D=0
M2952 868 115 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=52780 $D=0
M2953 869 115 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=57410 $D=0
M2954 870 115 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=62040 $D=0
M2955 871 115 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=66670 $D=0
M2956 202 116 872 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=52780 $D=0
M2957 203 116 873 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=57410 $D=0
M2958 204 116 874 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=62040 $D=0
M2959 205 116 875 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=66670 $D=0
M2960 876 117 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=52780 $D=0
M2961 877 117 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=57410 $D=0
M2962 878 117 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=62040 $D=0
M2963 879 117 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=66670 $D=0
M2964 880 872 280 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=52780 $D=0
M2965 881 873 281 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=57410 $D=0
M2966 882 874 282 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=62040 $D=0
M2967 883 875 283 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=66670 $D=0
M2968 202 880 1350 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=52780 $D=0
M2969 203 881 1351 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=57410 $D=0
M2970 204 882 1352 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=62040 $D=0
M2971 205 883 1353 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=66670 $D=0
M2972 884 1350 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=52780 $D=0
M2973 885 1351 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=57410 $D=0
M2974 886 1352 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=62040 $D=0
M2975 887 1353 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=66670 $D=0
M2976 880 116 884 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=52780 $D=0
M2977 881 116 885 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=57410 $D=0
M2978 882 116 886 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=62040 $D=0
M2979 883 116 887 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=66670 $D=0
M2980 884 876 300 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=52780 $D=0
M2981 885 877 301 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=57410 $D=0
M2982 886 878 302 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=62040 $D=0
M2983 887 879 303 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=66670 $D=0
M2984 308 888 884 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=52780 $D=0
M2985 309 889 885 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=57410 $D=0
M2986 310 890 886 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=62040 $D=0
M2987 311 891 887 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=66670 $D=0
M2988 888 118 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=52780 $D=0
M2989 889 118 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=57410 $D=0
M2990 890 118 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=62040 $D=0
M2991 891 118 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=66670 $D=0
M2992 202 119 892 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=52780 $D=0
M2993 203 119 893 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=57410 $D=0
M2994 204 119 894 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=62040 $D=0
M2995 205 119 895 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=66670 $D=0
M2996 896 120 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=52780 $D=0
M2997 897 120 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=57410 $D=0
M2998 898 120 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=62040 $D=0
M2999 899 120 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=66670 $D=0
M3000 900 892 280 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=52780 $D=0
M3001 901 893 281 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=57410 $D=0
M3002 902 894 282 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=62040 $D=0
M3003 903 895 283 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=66670 $D=0
M3004 202 900 1354 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=52780 $D=0
M3005 203 901 1355 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=57410 $D=0
M3006 204 902 1356 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=62040 $D=0
M3007 205 903 1357 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=66670 $D=0
M3008 904 1354 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=52780 $D=0
M3009 905 1355 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=57410 $D=0
M3010 906 1356 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=62040 $D=0
M3011 907 1357 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=66670 $D=0
M3012 900 119 904 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=52780 $D=0
M3013 901 119 905 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=57410 $D=0
M3014 902 119 906 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=62040 $D=0
M3015 903 119 907 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=66670 $D=0
M3016 904 896 300 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=52780 $D=0
M3017 905 897 301 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=57410 $D=0
M3018 906 898 302 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=62040 $D=0
M3019 907 899 303 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=66670 $D=0
M3020 308 908 904 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=52780 $D=0
M3021 309 909 905 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=57410 $D=0
M3022 310 910 906 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=62040 $D=0
M3023 311 911 907 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=66670 $D=0
M3024 908 121 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=52780 $D=0
M3025 909 121 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=57410 $D=0
M3026 910 121 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=62040 $D=0
M3027 911 121 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=66670 $D=0
M3028 202 122 912 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=52780 $D=0
M3029 203 122 913 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=57410 $D=0
M3030 204 122 914 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=62040 $D=0
M3031 205 122 915 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=66670 $D=0
M3032 916 123 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=52780 $D=0
M3033 917 123 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=57410 $D=0
M3034 918 123 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=62040 $D=0
M3035 919 123 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=66670 $D=0
M3036 8 916 300 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=52780 $D=0
M3037 9 917 301 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=57410 $D=0
M3038 10 918 302 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=62040 $D=0
M3039 11 919 303 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=66670 $D=0
M3040 308 912 8 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=52780 $D=0
M3041 309 913 9 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=57410 $D=0
M3042 310 914 10 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=62040 $D=0
M3043 311 915 11 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=66670 $D=0
M3044 202 924 920 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=52780 $D=0
M3045 203 925 921 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=57410 $D=0
M3046 204 926 922 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=62040 $D=0
M3047 205 927 923 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=66670 $D=0
M3048 924 124 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=52780 $D=0
M3049 925 124 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=57410 $D=0
M3050 926 124 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=62040 $D=0
M3051 927 124 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=66670 $D=0
M3052 1358 300 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=52780 $D=0
M3053 1359 301 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=57410 $D=0
M3054 1360 302 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=62040 $D=0
M3055 1361 303 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=66670 $D=0
M3056 928 924 1358 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=52780 $D=0
M3057 929 925 1359 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=57410 $D=0
M3058 930 926 1360 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=62040 $D=0
M3059 931 927 1361 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=66670 $D=0
M3060 202 928 932 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=52780 $D=0
M3061 203 929 933 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=57410 $D=0
M3062 204 930 934 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=62040 $D=0
M3063 205 931 935 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=66670 $D=0
M3064 1362 932 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=52780 $D=0
M3065 1363 933 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=57410 $D=0
M3066 1364 934 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=62040 $D=0
M3067 1365 935 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=66670 $D=0
M3068 928 920 1362 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=52780 $D=0
M3069 929 921 1363 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=57410 $D=0
M3070 930 922 1364 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=62040 $D=0
M3071 931 923 1365 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=66670 $D=0
M3072 202 940 936 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=52780 $D=0
M3073 203 941 937 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=57410 $D=0
M3074 204 942 938 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=62040 $D=0
M3075 205 943 939 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=66670 $D=0
M3076 940 124 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=52780 $D=0
M3077 941 124 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=57410 $D=0
M3078 942 124 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=62040 $D=0
M3079 943 124 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=66670 $D=0
M3080 1366 308 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=52780 $D=0
M3081 1367 309 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=57410 $D=0
M3082 1368 310 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=62040 $D=0
M3083 1369 311 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=66670 $D=0
M3084 944 940 1366 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=52780 $D=0
M3085 945 941 1367 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=57410 $D=0
M3086 946 942 1368 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=62040 $D=0
M3087 947 943 1369 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=66670 $D=0
M3088 202 944 125 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=52780 $D=0
M3089 203 945 126 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=57410 $D=0
M3090 204 946 127 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=62040 $D=0
M3091 205 947 128 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=66670 $D=0
M3092 1370 125 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=52780 $D=0
M3093 1371 126 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=57410 $D=0
M3094 1372 127 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=62040 $D=0
M3095 1373 128 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=66670 $D=0
M3096 944 936 1370 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=52780 $D=0
M3097 945 937 1371 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=57410 $D=0
M3098 946 938 1372 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=62040 $D=0
M3099 947 939 1373 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=66670 $D=0
M3100 948 129 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=52780 $D=0
M3101 949 129 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=57410 $D=0
M3102 950 129 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=62040 $D=0
M3103 951 129 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=66670 $D=0
M3104 952 129 932 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=52780 $D=0
M3105 953 129 933 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=57410 $D=0
M3106 954 129 934 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=62040 $D=0
M3107 955 129 935 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=66670 $D=0
M3108 130 948 952 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=52780 $D=0
M3109 131 949 953 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=57410 $D=0
M3110 132 950 954 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=62040 $D=0
M3111 133 951 955 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=66670 $D=0
M3112 956 134 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=52780 $D=0
M3113 957 134 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=57410 $D=0
M3114 958 134 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=62040 $D=0
M3115 959 134 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=66670 $D=0
M3116 960 134 125 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=52780 $D=0
M3117 961 134 126 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=57410 $D=0
M3118 962 134 127 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=62040 $D=0
M3119 963 134 128 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=66670 $D=0
M3120 1374 956 960 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=52780 $D=0
M3121 1375 957 961 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=57410 $D=0
M3122 1376 958 962 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=62040 $D=0
M3123 1377 959 963 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=66670 $D=0
M3124 202 125 1374 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=52780 $D=0
M3125 203 126 1375 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=57410 $D=0
M3126 204 127 1376 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=62040 $D=0
M3127 205 128 1377 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=66670 $D=0
M3128 964 135 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=52780 $D=0
M3129 965 135 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=57410 $D=0
M3130 966 135 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=62040 $D=0
M3131 967 135 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=66670 $D=0
M3132 968 135 960 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=52780 $D=0
M3133 969 135 961 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=57410 $D=0
M3134 970 135 962 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=62040 $D=0
M3135 971 135 963 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=66670 $D=0
M3136 15 964 968 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=52780 $D=0
M3137 16 965 969 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=57410 $D=0
M3138 17 966 970 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=62040 $D=0
M3139 18 967 971 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=66670 $D=0
M3140 975 972 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=52780 $D=0
M3141 976 973 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=57410 $D=0
M3142 977 974 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=62040 $D=0
M3143 978 136 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=66670 $D=0
M3144 202 983 979 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=52780 $D=0
M3145 203 984 980 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=57410 $D=0
M3146 204 985 981 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=62040 $D=0
M3147 205 986 982 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=66670 $D=0
M3148 987 952 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=52780 $D=0
M3149 988 953 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=57410 $D=0
M3150 989 954 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=62040 $D=0
M3151 990 955 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=66670 $D=0
M3152 983 952 972 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=52780 $D=0
M3153 984 953 973 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=57410 $D=0
M3154 985 954 974 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=62040 $D=0
M3155 986 955 136 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=66670 $D=0
M3156 975 987 983 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=52780 $D=0
M3157 976 988 984 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=57410 $D=0
M3158 977 989 985 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=62040 $D=0
M3159 978 990 986 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=66670 $D=0
M3160 991 979 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=52780 $D=0
M3161 992 980 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=57410 $D=0
M3162 993 981 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=62040 $D=0
M3163 994 982 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=66670 $D=0
M3164 137 979 968 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=52780 $D=0
M3165 972 980 969 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=57410 $D=0
M3166 973 981 970 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=62040 $D=0
M3167 974 982 971 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=66670 $D=0
M3168 952 991 137 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=52780 $D=0
M3169 953 992 972 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=57410 $D=0
M3170 954 993 973 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=62040 $D=0
M3171 955 994 974 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=66670 $D=0
M3172 995 137 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=52780 $D=0
M3173 996 972 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=57410 $D=0
M3174 997 973 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=62040 $D=0
M3175 998 974 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=66670 $D=0
M3176 999 979 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=52780 $D=0
M3177 1000 980 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=57410 $D=0
M3178 1001 981 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=62040 $D=0
M3179 1002 982 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=66670 $D=0
M3180 1003 979 995 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=52780 $D=0
M3181 1004 980 996 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=57410 $D=0
M3182 1005 981 997 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=62040 $D=0
M3183 1006 982 998 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=66670 $D=0
M3184 968 999 1003 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=52780 $D=0
M3185 969 1000 1004 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=57410 $D=0
M3186 970 1001 1005 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=62040 $D=0
M3187 971 1002 1006 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=66670 $D=0
M3188 1410 952 202 202 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=52420 $D=0
M3189 1411 953 203 203 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=57050 $D=0
M3190 1412 954 204 204 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=61680 $D=0
M3191 1413 955 205 205 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=66310 $D=0
M3192 1007 968 1410 202 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=52420 $D=0
M3193 1008 969 1411 203 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=57050 $D=0
M3194 1009 970 1412 204 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=61680 $D=0
M3195 1010 971 1413 205 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=66310 $D=0
M3196 1011 1003 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=52780 $D=0
M3197 1012 1004 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=57410 $D=0
M3198 1013 1005 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=62040 $D=0
M3199 1014 1006 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=66670 $D=0
M3200 1015 952 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=52780 $D=0
M3201 1016 953 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=57410 $D=0
M3202 1017 954 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=62040 $D=0
M3203 1018 955 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=66670 $D=0
M3204 202 968 1015 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=52780 $D=0
M3205 203 969 1016 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=57410 $D=0
M3206 204 970 1017 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=62040 $D=0
M3207 205 971 1018 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=66670 $D=0
M3208 1019 952 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=52780 $D=0
M3209 1020 953 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=57410 $D=0
M3210 1021 954 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=62040 $D=0
M3211 1022 955 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=66670 $D=0
M3212 202 968 1019 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=52780 $D=0
M3213 203 969 1020 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=57410 $D=0
M3214 204 970 1021 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=62040 $D=0
M3215 205 971 1022 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=66670 $D=0
M3216 1414 952 202 202 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=52600 $D=0
M3217 1415 953 203 203 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=57230 $D=0
M3218 1416 954 204 204 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=61860 $D=0
M3219 1417 955 205 205 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=66490 $D=0
M3220 1027 968 1414 202 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=52600 $D=0
M3221 1028 969 1415 203 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=57230 $D=0
M3222 1029 970 1416 204 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=61860 $D=0
M3223 1030 971 1417 205 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=66490 $D=0
M3224 202 1019 1027 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=52780 $D=0
M3225 203 1020 1028 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=57410 $D=0
M3226 204 1021 1029 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=62040 $D=0
M3227 205 1022 1030 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=66670 $D=0
M3228 1031 144 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=52780 $D=0
M3229 1032 144 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=57410 $D=0
M3230 1033 144 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=62040 $D=0
M3231 1034 144 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=66670 $D=0
M3232 1035 144 1007 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=52780 $D=0
M3233 1036 144 1008 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=57410 $D=0
M3234 1037 144 1009 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=62040 $D=0
M3235 1038 144 1010 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=66670 $D=0
M3236 1015 1031 1035 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=52780 $D=0
M3237 1016 1032 1036 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=57410 $D=0
M3238 1017 1033 1037 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=62040 $D=0
M3239 1018 1034 1038 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=66670 $D=0
M3240 1039 144 1011 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=52780 $D=0
M3241 1040 144 1012 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=57410 $D=0
M3242 1041 144 1013 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=62040 $D=0
M3243 1042 144 1014 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=66670 $D=0
M3244 1027 1031 1039 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=52780 $D=0
M3245 1028 1032 1040 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=57410 $D=0
M3246 1029 1033 1041 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=62040 $D=0
M3247 1030 1034 1042 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=66670 $D=0
M3248 1043 145 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=52780 $D=0
M3249 1044 145 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=57410 $D=0
M3250 1045 145 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=62040 $D=0
M3251 1046 145 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=66670 $D=0
M3252 1047 145 1039 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=52780 $D=0
M3253 1048 145 1040 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=57410 $D=0
M3254 1049 145 1041 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=62040 $D=0
M3255 1050 145 1042 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=66670 $D=0
M3256 1035 1043 1047 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=52780 $D=0
M3257 1036 1044 1048 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=57410 $D=0
M3258 1037 1045 1049 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=62040 $D=0
M3259 1038 1046 1050 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=66670 $D=0
M3260 19 1047 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=52780 $D=0
M3261 20 1048 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=57410 $D=0
M3262 21 1049 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=62040 $D=0
M3263 22 1050 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=66670 $D=0
M3264 1051 146 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=52780 $D=0
M3265 1052 146 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=57410 $D=0
M3266 1053 146 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=62040 $D=0
M3267 1054 146 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=66670 $D=0
M3268 1055 146 147 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=52780 $D=0
M3269 1056 146 148 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=57410 $D=0
M3270 1057 146 149 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=62040 $D=0
M3271 1058 146 150 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=66670 $D=0
M3272 151 1051 1055 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=52780 $D=0
M3273 152 1052 1056 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=57410 $D=0
M3274 147 1053 1057 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=62040 $D=0
M3275 148 1054 1058 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=66670 $D=0
M3276 1059 146 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=52780 $D=0
M3277 1060 146 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=57410 $D=0
M3278 1061 146 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=62040 $D=0
M3279 1062 146 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=66670 $D=0
M3280 1064 146 153 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=52780 $D=0
M3281 1065 146 155 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=57410 $D=0
M3282 1066 146 156 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=62040 $D=0
M3283 1067 146 158 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=66670 $D=0
M3284 159 1059 1064 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=52780 $D=0
M3285 154 1060 1065 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=57410 $D=0
M3286 160 1061 1066 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=62040 $D=0
M3287 157 1062 1067 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=66670 $D=0
M3288 1068 146 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=52780 $D=0
M3289 1069 146 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=57410 $D=0
M3290 1070 146 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=62040 $D=0
M3291 1071 146 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=66670 $D=0
M3292 1072 146 138 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=52780 $D=0
M3293 1073 146 143 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=57410 $D=0
M3294 1074 146 141 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=62040 $D=0
M3295 1075 146 161 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=66670 $D=0
M3296 162 1068 1072 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=52780 $D=0
M3297 163 1069 1073 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=57410 $D=0
M3298 164 1070 1074 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=62040 $D=0
M3299 165 1071 1075 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=66670 $D=0
M3300 1076 146 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=52780 $D=0
M3301 1077 146 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=57410 $D=0
M3302 1078 146 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=62040 $D=0
M3303 1079 146 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=66670 $D=0
M3304 1080 146 166 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=52780 $D=0
M3305 1081 146 167 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=57410 $D=0
M3306 1082 146 168 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=62040 $D=0
M3307 1083 146 169 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=66670 $D=0
M3308 170 1076 1080 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=52780 $D=0
M3309 171 1077 1081 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=57410 $D=0
M3310 172 1078 1082 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=62040 $D=0
M3311 173 1079 1083 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=66670 $D=0
M3312 1084 146 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=52780 $D=0
M3313 1085 146 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=57410 $D=0
M3314 1086 146 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=62040 $D=0
M3315 1087 146 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=66670 $D=0
M3316 1088 146 174 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=52780 $D=0
M3317 1089 146 175 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=57410 $D=0
M3318 1090 146 176 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=62040 $D=0
M3319 1091 146 177 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=66670 $D=0
M3320 178 1084 1088 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=52780 $D=0
M3321 178 1085 1089 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=57410 $D=0
M3322 178 1086 1090 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=62040 $D=0
M3323 178 1087 1091 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=66670 $D=0
M3324 202 952 1390 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=52780 $D=0
M3325 203 953 1391 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=57410 $D=0
M3326 204 954 1392 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=62040 $D=0
M3327 205 955 1393 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=66670 $D=0
M3328 152 1390 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=52780 $D=0
M3329 147 1391 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=57410 $D=0
M3330 148 1392 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=62040 $D=0
M3331 149 1393 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=66670 $D=0
M3332 1092 179 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=52780 $D=0
M3333 1093 179 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=57410 $D=0
M3334 1094 179 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=62040 $D=0
M3335 1095 179 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=66670 $D=0
M3336 160 179 152 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=52780 $D=0
M3337 157 179 147 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=57410 $D=0
M3338 153 179 148 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=62040 $D=0
M3339 155 179 149 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=66670 $D=0
M3340 1055 1092 160 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=52780 $D=0
M3341 1056 1093 157 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=57410 $D=0
M3342 1057 1094 153 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=62040 $D=0
M3343 1058 1095 155 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=66670 $D=0
M3344 1096 180 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=52780 $D=0
M3345 1097 180 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=57410 $D=0
M3346 1098 180 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=62040 $D=0
M3347 1099 180 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=66670 $D=0
M3348 181 180 160 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=52780 $D=0
M3349 142 180 157 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=57410 $D=0
M3350 140 180 153 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=62040 $D=0
M3351 139 180 155 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=66670 $D=0
M3352 1064 1096 181 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=52780 $D=0
M3353 1065 1097 142 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=57410 $D=0
M3354 1066 1098 140 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=62040 $D=0
M3355 1067 1099 139 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=66670 $D=0
M3356 1100 182 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=52780 $D=0
M3357 1101 182 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=57410 $D=0
M3358 1102 182 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=62040 $D=0
M3359 1103 182 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=66670 $D=0
M3360 183 182 181 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=52780 $D=0
M3361 184 182 142 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=57410 $D=0
M3362 185 182 140 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=62040 $D=0
M3363 186 182 139 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=66670 $D=0
M3364 1072 1100 183 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=52780 $D=0
M3365 1073 1101 184 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=57410 $D=0
M3366 1074 1102 185 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=62040 $D=0
M3367 1075 1103 186 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=66670 $D=0
M3368 1104 187 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=52780 $D=0
M3369 1105 187 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=57410 $D=0
M3370 1106 187 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=62040 $D=0
M3371 1107 187 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=66670 $D=0
M3372 188 187 183 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=52780 $D=0
M3373 189 187 184 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=57410 $D=0
M3374 190 187 185 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=62040 $D=0
M3375 191 187 186 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=66670 $D=0
M3376 1080 1104 188 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=52780 $D=0
M3377 1081 1105 189 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=57410 $D=0
M3378 1082 1106 190 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=62040 $D=0
M3379 1083 1107 191 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=66670 $D=0
M3380 1108 192 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=52780 $D=0
M3381 1109 192 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=57410 $D=0
M3382 1110 192 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=62040 $D=0
M3383 1111 192 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=66670 $D=0
M3384 23 192 188 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=52780 $D=0
M3385 24 192 189 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=57410 $D=0
M3386 25 192 190 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=62040 $D=0
M3387 26 192 191 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=66670 $D=0
M3388 1088 1108 23 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=52780 $D=0
M3389 1089 1109 24 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=57410 $D=0
M3390 1090 1110 25 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=62040 $D=0
M3391 1091 1111 26 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=66670 $D=0
M3392 1112 193 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=52780 $D=0
M3393 1113 193 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=57410 $D=0
M3394 1114 193 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=62040 $D=0
M3395 1115 193 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=66670 $D=0
M3396 1116 193 125 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=52780 $D=0
M3397 1117 193 126 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=57410 $D=0
M3398 1118 193 127 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=62040 $D=0
M3399 1119 193 128 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=66670 $D=0
M3400 15 1112 1116 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=52780 $D=0
M3401 16 1113 1117 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=57410 $D=0
M3402 17 1114 1118 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=62040 $D=0
M3403 18 1115 1119 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=66670 $D=0
M3404 1120 932 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=52780 $D=0
M3405 1121 933 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=57410 $D=0
M3406 1122 934 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=62040 $D=0
M3407 1123 935 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=66670 $D=0
M3408 202 1116 1120 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=52780 $D=0
M3409 203 1117 1121 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=57410 $D=0
M3410 204 1118 1122 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=62040 $D=0
M3411 205 1119 1123 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=66670 $D=0
M3412 1418 932 202 202 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=52600 $D=0
M3413 1419 933 203 203 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=57230 $D=0
M3414 1420 934 204 204 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=61860 $D=0
M3415 1421 935 205 205 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=66490 $D=0
M3416 1128 1116 1418 202 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=52600 $D=0
M3417 1129 1117 1419 203 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=57230 $D=0
M3418 1130 1118 1420 204 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=61860 $D=0
M3419 1131 1119 1421 205 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=66490 $D=0
M3420 202 1120 1128 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=52780 $D=0
M3421 203 1121 1129 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=57410 $D=0
M3422 204 1122 1130 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=62040 $D=0
M3423 205 1123 1131 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=66670 $D=0
M3424 1394 194 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=52780 $D=0
M3425 1395 1132 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=57410 $D=0
M3426 1396 1133 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=62040 $D=0
M3427 1397 1134 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=66670 $D=0
M3428 202 1128 1394 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=52780 $D=0
M3429 203 1129 1395 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=57410 $D=0
M3430 204 1130 1396 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=62040 $D=0
M3431 205 1131 1397 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=66670 $D=0
M3432 1132 1394 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=52780 $D=0
M3433 1135 1395 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=57410 $D=0
M3434 1134 1396 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=62040 $D=0
M3435 195 1397 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=66670 $D=0
M3436 1422 932 202 202 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=52420 $D=0
M3437 1423 933 203 203 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=57050 $D=0
M3438 1424 934 204 204 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=61680 $D=0
M3439 1425 935 205 205 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=66310 $D=0
M3440 1136 1140 1422 202 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=52420 $D=0
M3441 1137 1141 1423 203 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=57050 $D=0
M3442 1138 1142 1424 204 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=61680 $D=0
M3443 1139 1143 1425 205 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=66310 $D=0
M3444 1140 1116 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=52780 $D=0
M3445 1141 1117 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=57410 $D=0
M3446 1142 1118 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=62040 $D=0
M3447 1143 1119 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=66670 $D=0
M3448 1144 1136 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=52780 $D=0
M3449 1145 1137 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=57410 $D=0
M3450 1146 1138 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=62040 $D=0
M3451 1147 1139 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=66670 $D=0
M3452 202 194 1144 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=52780 $D=0
M3453 203 1132 1145 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=57410 $D=0
M3454 204 1133 1146 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=62040 $D=0
M3455 205 1134 1147 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=66670 $D=0
M3456 1151 196 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=52780 $D=0
M3457 1152 1148 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=57410 $D=0
M3458 1153 1149 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=62040 $D=0
M3459 1154 1150 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=66670 $D=0
M3460 1148 1144 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=52780 $D=0
M3461 1149 1145 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=57410 $D=0
M3462 1150 1146 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=62040 $D=0
M3463 197 1147 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=66670 $D=0
M3464 202 1151 1148 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=52780 $D=0
M3465 203 1152 1149 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=57410 $D=0
M3466 204 1153 1150 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=62040 $D=0
M3467 205 1154 197 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=66670 $D=0
M3468 1158 1155 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=52780 $D=0
M3469 1159 1156 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=57410 $D=0
M3470 1160 1157 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=62040 $D=0
M3471 1161 198 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=66670 $D=0
M3472 202 1166 1162 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=52780 $D=0
M3473 203 1167 1163 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=57410 $D=0
M3474 204 1168 1164 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=62040 $D=0
M3475 205 1169 1165 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=66670 $D=0
M3476 1170 130 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=52780 $D=0
M3477 1171 131 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=57410 $D=0
M3478 1172 132 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=62040 $D=0
M3479 1173 133 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=66670 $D=0
M3480 1166 130 1155 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=52780 $D=0
M3481 1167 131 1156 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=57410 $D=0
M3482 1168 132 1157 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=62040 $D=0
M3483 1169 133 198 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=66670 $D=0
M3484 1158 1170 1166 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=52780 $D=0
M3485 1159 1171 1167 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=57410 $D=0
M3486 1160 1172 1168 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=62040 $D=0
M3487 1161 1173 1169 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=66670 $D=0
M3488 1174 1162 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=52780 $D=0
M3489 1175 1163 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=57410 $D=0
M3490 1176 1164 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=62040 $D=0
M3491 1177 1165 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=66670 $D=0
M3492 199 1162 8 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=52780 $D=0
M3493 1155 1163 9 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=57410 $D=0
M3494 1156 1164 10 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=62040 $D=0
M3495 1157 1165 11 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=66670 $D=0
M3496 130 1174 199 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=52780 $D=0
M3497 131 1175 1155 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=57410 $D=0
M3498 132 1176 1156 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=62040 $D=0
M3499 133 1177 1157 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=66670 $D=0
M3500 1178 199 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=52780 $D=0
M3501 1179 1155 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=57410 $D=0
M3502 1180 1156 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=62040 $D=0
M3503 1181 1157 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=66670 $D=0
M3504 1182 1162 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=52780 $D=0
M3505 1183 1163 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=57410 $D=0
M3506 1184 1164 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=62040 $D=0
M3507 1185 1165 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=66670 $D=0
M3508 256 1162 1178 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=52780 $D=0
M3509 257 1163 1179 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=57410 $D=0
M3510 258 1164 1180 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=62040 $D=0
M3511 259 1165 1181 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=66670 $D=0
M3512 8 1182 256 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=52780 $D=0
M3513 9 1183 257 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=57410 $D=0
M3514 10 1184 258 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=62040 $D=0
M3515 11 1185 259 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=66670 $D=0
M3516 1186 200 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=52780 $D=0
M3517 1187 200 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=57410 $D=0
M3518 1188 200 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=62040 $D=0
M3519 1189 200 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=66670 $D=0
M3520 1190 200 256 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=52780 $D=0
M3521 1191 200 257 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=57410 $D=0
M3522 1192 200 258 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=62040 $D=0
M3523 1193 200 259 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=66670 $D=0
M3524 19 1186 1190 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=52780 $D=0
M3525 20 1187 1191 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=57410 $D=0
M3526 21 1188 1192 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=62040 $D=0
M3527 22 1189 1193 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=66670 $D=0
M3528 1194 201 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=52780 $D=0
M3529 1195 201 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=57410 $D=0
M3530 1196 201 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=62040 $D=0
M3531 1197 201 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=66670 $D=0
M3532 201 201 1190 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=52780 $D=0
M3533 201 201 1191 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=57410 $D=0
M3534 201 201 1192 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=62040 $D=0
M3535 201 201 1193 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=66670 $D=0
M3536 8 1194 201 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=52780 $D=0
M3537 9 1195 201 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=57410 $D=0
M3538 10 1196 201 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=62040 $D=0
M3539 11 1197 201 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=66670 $D=0
M3540 1198 124 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=52780 $D=0
M3541 1199 124 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=57410 $D=0
M3542 1200 124 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=62040 $D=0
M3543 1201 124 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=66670 $D=0
M3544 202 1198 1202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=52780 $D=0
M3545 203 1199 1203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=57410 $D=0
M3546 204 1200 1204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=62040 $D=0
M3547 205 1201 1205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=66670 $D=0
M3548 1206 124 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=52780 $D=0
M3549 1207 124 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=57410 $D=0
M3550 1208 124 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=62040 $D=0
M3551 1209 124 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=66670 $D=0
M3552 1210 1202 201 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=52780 $D=0
M3553 1211 1203 201 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=57410 $D=0
M3554 1212 1204 201 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=62040 $D=0
M3555 1213 1205 201 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=66670 $D=0
M3556 202 1210 1398 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=52780 $D=0
M3557 203 1211 1399 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=57410 $D=0
M3558 204 1212 1400 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=62040 $D=0
M3559 205 1213 1401 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=66670 $D=0
M3560 1214 1398 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=52780 $D=0
M3561 1215 1399 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=57410 $D=0
M3562 1216 1400 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=62040 $D=0
M3563 1217 1401 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=66670 $D=0
M3564 1210 1198 1214 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=52780 $D=0
M3565 1211 1199 1215 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=57410 $D=0
M3566 1212 1200 1216 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=62040 $D=0
M3567 1213 1201 1217 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=66670 $D=0
M3568 1218 1206 1214 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=52780 $D=0
M3569 1219 1207 1215 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=57410 $D=0
M3570 1220 1208 1216 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=62040 $D=0
M3571 1221 1209 1217 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=66670 $D=0
M3572 202 1226 1222 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=52780 $D=0
M3573 203 1227 1223 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=57410 $D=0
M3574 204 1228 1224 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=62040 $D=0
M3575 205 1229 1225 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=66670 $D=0
M3576 1226 124 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=52780 $D=0
M3577 1227 124 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=57410 $D=0
M3578 1228 124 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=62040 $D=0
M3579 1229 124 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=66670 $D=0
M3580 1402 1218 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=52780 $D=0
M3581 1403 1219 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=57410 $D=0
M3582 1404 1220 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=62040 $D=0
M3583 1405 1221 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=66670 $D=0
M3584 1230 1226 1402 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=52780 $D=0
M3585 1231 1227 1403 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=57410 $D=0
M3586 1232 1228 1404 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=62040 $D=0
M3587 1233 1229 1405 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=66670 $D=0
M3588 202 1230 130 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=52780 $D=0
M3589 203 1231 131 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=57410 $D=0
M3590 204 1232 132 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=62040 $D=0
M3591 205 1233 133 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=66670 $D=0
M3592 1406 130 202 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=52780 $D=0
M3593 1407 131 203 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=57410 $D=0
M3594 1408 132 204 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=62040 $D=0
M3595 1409 133 205 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=66670 $D=0
M3596 1230 1222 1406 202 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=52780 $D=0
M3597 1231 1223 1407 203 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=57410 $D=0
M3598 1232 1224 1408 204 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=62040 $D=0
M3599 1233 1225 1409 205 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=66670 $D=0
.ENDS
***************************************
.SUBCKT ICV_37 1 2 3 4 5 6 7 9 10 11 12 13 14 15 16 17 18 19 20 21
+ 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41
+ 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61
+ 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81
+ 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101
+ 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121
+ 122 123 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141 142
+ 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162
+ 163 164 165 166 167 168 169
** N=797 EP=167 IP=1514 FDC=1800
M0 175 1 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=42270 $D=1
M1 176 1 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=46900 $D=1
M2 177 175 2 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=42270 $D=1
M3 178 176 3 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=46900 $D=1
M4 6 1 177 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=42270 $D=1
M5 7 1 178 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=46900 $D=1
M6 179 175 4 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=42270 $D=1
M7 180 176 4 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=46900 $D=1
M8 5 1 179 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=42270 $D=1
M9 5 1 180 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=46900 $D=1
M10 181 175 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=42270 $D=1
M11 182 176 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=46900 $D=1
M12 6 1 181 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=42270 $D=1
M13 7 1 182 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=46900 $D=1
M14 185 183 181 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=42270 $D=1
M15 186 184 182 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=46900 $D=1
M16 183 9 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=42270 $D=1
M17 184 9 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=46900 $D=1
M18 187 183 179 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=42270 $D=1
M19 188 184 180 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=46900 $D=1
M20 177 9 187 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=42270 $D=1
M21 178 9 188 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=46900 $D=1
M22 189 10 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=42270 $D=1
M23 190 10 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=46900 $D=1
M24 191 189 187 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=42270 $D=1
M25 192 190 188 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=46900 $D=1
M26 185 10 191 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=42270 $D=1
M27 186 10 192 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=46900 $D=1
M28 193 11 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=42270 $D=1
M29 194 11 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=46900 $D=1
M30 195 193 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=42270 $D=1
M31 196 194 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=46900 $D=1
M32 12 11 195 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=42270 $D=1
M33 13 11 196 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=46900 $D=1
M34 197 193 14 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=42270 $D=1
M35 198 194 15 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=46900 $D=1
M36 16 11 197 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=42270 $D=1
M37 17 11 198 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=46900 $D=1
M38 201 193 199 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=42270 $D=1
M39 202 194 200 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=46900 $D=1
M40 191 11 201 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=42270 $D=1
M41 192 11 202 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=46900 $D=1
M42 205 203 201 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=42270 $D=1
M43 206 204 202 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=46900 $D=1
M44 203 18 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=42270 $D=1
M45 204 18 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=46900 $D=1
M46 207 203 197 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=42270 $D=1
M47 208 204 198 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=46900 $D=1
M48 195 18 207 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=42270 $D=1
M49 196 18 208 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=46900 $D=1
M50 209 19 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=42270 $D=1
M51 210 19 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=46900 $D=1
M52 211 209 207 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=42270 $D=1
M53 212 210 208 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=46900 $D=1
M54 205 19 211 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=42270 $D=1
M55 206 19 212 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=46900 $D=1
M56 6 20 213 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=42270 $D=1
M57 7 20 214 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=46900 $D=1
M58 215 21 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=42270 $D=1
M59 216 21 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=46900 $D=1
M60 217 20 211 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=42270 $D=1
M61 218 20 212 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=46900 $D=1
M62 6 217 688 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=42270 $D=1
M63 7 218 689 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=46900 $D=1
M64 219 688 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=42270 $D=1
M65 220 689 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=46900 $D=1
M66 217 213 219 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=42270 $D=1
M67 218 214 220 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=46900 $D=1
M68 219 21 221 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=42270 $D=1
M69 220 21 222 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=46900 $D=1
M70 225 22 219 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=42270 $D=1
M71 226 22 220 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=46900 $D=1
M72 223 22 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=42270 $D=1
M73 224 22 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=46900 $D=1
M74 6 23 227 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=42270 $D=1
M75 7 23 228 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=46900 $D=1
M76 229 24 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=42270 $D=1
M77 230 24 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=46900 $D=1
M78 231 23 211 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=42270 $D=1
M79 232 23 212 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=46900 $D=1
M80 6 231 690 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=42270 $D=1
M81 7 232 691 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=46900 $D=1
M82 233 690 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=42270 $D=1
M83 234 691 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=46900 $D=1
M84 231 227 233 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=42270 $D=1
M85 232 228 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=46900 $D=1
M86 233 24 221 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=42270 $D=1
M87 234 24 222 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=46900 $D=1
M88 225 25 233 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=42270 $D=1
M89 226 25 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=46900 $D=1
M90 235 25 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=42270 $D=1
M91 236 25 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=46900 $D=1
M92 6 26 237 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=42270 $D=1
M93 7 26 238 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=46900 $D=1
M94 239 27 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=42270 $D=1
M95 240 27 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=46900 $D=1
M96 241 26 211 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=42270 $D=1
M97 242 26 212 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=46900 $D=1
M98 6 241 692 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=42270 $D=1
M99 7 242 693 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=46900 $D=1
M100 243 692 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=42270 $D=1
M101 244 693 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=46900 $D=1
M102 241 237 243 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=42270 $D=1
M103 242 238 244 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=46900 $D=1
M104 243 27 221 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=42270 $D=1
M105 244 27 222 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=46900 $D=1
M106 225 28 243 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=42270 $D=1
M107 226 28 244 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=46900 $D=1
M108 245 28 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=42270 $D=1
M109 246 28 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=46900 $D=1
M110 6 29 247 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=42270 $D=1
M111 7 29 248 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=46900 $D=1
M112 249 30 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=42270 $D=1
M113 250 30 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=46900 $D=1
M114 251 29 211 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=42270 $D=1
M115 252 29 212 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=46900 $D=1
M116 6 251 694 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=42270 $D=1
M117 7 252 695 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=46900 $D=1
M118 253 694 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=42270 $D=1
M119 254 695 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=46900 $D=1
M120 251 247 253 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=42270 $D=1
M121 252 248 254 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=46900 $D=1
M122 253 30 221 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=42270 $D=1
M123 254 30 222 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=46900 $D=1
M124 225 31 253 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=42270 $D=1
M125 226 31 254 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=46900 $D=1
M126 255 31 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=42270 $D=1
M127 256 31 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=46900 $D=1
M128 6 32 257 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=42270 $D=1
M129 7 32 258 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=46900 $D=1
M130 259 33 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=42270 $D=1
M131 260 33 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=46900 $D=1
M132 261 32 211 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=42270 $D=1
M133 262 32 212 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=46900 $D=1
M134 6 261 696 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=42270 $D=1
M135 7 262 697 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=46900 $D=1
M136 263 696 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=42270 $D=1
M137 264 697 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=46900 $D=1
M138 261 257 263 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=42270 $D=1
M139 262 258 264 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=46900 $D=1
M140 263 33 221 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=42270 $D=1
M141 264 33 222 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=46900 $D=1
M142 225 34 263 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=42270 $D=1
M143 226 34 264 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=46900 $D=1
M144 265 34 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=42270 $D=1
M145 266 34 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=46900 $D=1
M146 6 35 267 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=42270 $D=1
M147 7 35 268 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=46900 $D=1
M148 269 36 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=42270 $D=1
M149 270 36 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=46900 $D=1
M150 271 35 211 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=42270 $D=1
M151 272 35 212 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=46900 $D=1
M152 6 271 698 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=42270 $D=1
M153 7 272 699 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=46900 $D=1
M154 273 698 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=42270 $D=1
M155 274 699 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=46900 $D=1
M156 271 267 273 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=42270 $D=1
M157 272 268 274 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=46900 $D=1
M158 273 36 221 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=42270 $D=1
M159 274 36 222 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=46900 $D=1
M160 225 37 273 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=42270 $D=1
M161 226 37 274 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=46900 $D=1
M162 275 37 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=42270 $D=1
M163 276 37 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=46900 $D=1
M164 6 38 277 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=42270 $D=1
M165 7 38 278 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=46900 $D=1
M166 279 39 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=42270 $D=1
M167 280 39 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=46900 $D=1
M168 281 38 211 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=42270 $D=1
M169 282 38 212 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=46900 $D=1
M170 6 281 700 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=42270 $D=1
M171 7 282 701 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=46900 $D=1
M172 283 700 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=42270 $D=1
M173 284 701 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=46900 $D=1
M174 281 277 283 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=42270 $D=1
M175 282 278 284 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=46900 $D=1
M176 283 39 221 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=42270 $D=1
M177 284 39 222 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=46900 $D=1
M178 225 40 283 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=42270 $D=1
M179 226 40 284 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=46900 $D=1
M180 285 40 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=42270 $D=1
M181 286 40 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=46900 $D=1
M182 6 41 287 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=42270 $D=1
M183 7 41 288 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=46900 $D=1
M184 289 42 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=42270 $D=1
M185 290 42 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=46900 $D=1
M186 291 41 211 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=42270 $D=1
M187 292 41 212 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=46900 $D=1
M188 6 291 702 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=42270 $D=1
M189 7 292 703 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=46900 $D=1
M190 293 702 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=42270 $D=1
M191 294 703 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=46900 $D=1
M192 291 287 293 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=42270 $D=1
M193 292 288 294 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=46900 $D=1
M194 293 42 221 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=42270 $D=1
M195 294 42 222 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=46900 $D=1
M196 225 43 293 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=42270 $D=1
M197 226 43 294 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=46900 $D=1
M198 295 43 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=42270 $D=1
M199 296 43 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=46900 $D=1
M200 6 44 297 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=42270 $D=1
M201 7 44 298 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=46900 $D=1
M202 299 45 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=42270 $D=1
M203 300 45 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=46900 $D=1
M204 301 44 211 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=42270 $D=1
M205 302 44 212 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=46900 $D=1
M206 6 301 704 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=42270 $D=1
M207 7 302 705 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=46900 $D=1
M208 303 704 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=42270 $D=1
M209 304 705 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=46900 $D=1
M210 301 297 303 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=42270 $D=1
M211 302 298 304 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=46900 $D=1
M212 303 45 221 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=42270 $D=1
M213 304 45 222 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=46900 $D=1
M214 225 46 303 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=42270 $D=1
M215 226 46 304 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=46900 $D=1
M216 305 46 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=42270 $D=1
M217 306 46 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=46900 $D=1
M218 6 47 307 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=42270 $D=1
M219 7 47 308 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=46900 $D=1
M220 309 48 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=42270 $D=1
M221 310 48 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=46900 $D=1
M222 311 47 211 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=42270 $D=1
M223 312 47 212 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=46900 $D=1
M224 6 311 706 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=42270 $D=1
M225 7 312 707 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=46900 $D=1
M226 313 706 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=42270 $D=1
M227 314 707 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=46900 $D=1
M228 311 307 313 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=42270 $D=1
M229 312 308 314 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=46900 $D=1
M230 313 48 221 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=42270 $D=1
M231 314 48 222 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=46900 $D=1
M232 225 49 313 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=42270 $D=1
M233 226 49 314 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=46900 $D=1
M234 315 49 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=42270 $D=1
M235 316 49 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=46900 $D=1
M236 6 50 317 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=42270 $D=1
M237 7 50 318 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=46900 $D=1
M238 319 51 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=42270 $D=1
M239 320 51 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=46900 $D=1
M240 321 50 211 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=42270 $D=1
M241 322 50 212 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=46900 $D=1
M242 6 321 708 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=42270 $D=1
M243 7 322 709 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=46900 $D=1
M244 323 708 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=42270 $D=1
M245 324 709 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=46900 $D=1
M246 321 317 323 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=42270 $D=1
M247 322 318 324 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=46900 $D=1
M248 323 51 221 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=42270 $D=1
M249 324 51 222 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=46900 $D=1
M250 225 52 323 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=42270 $D=1
M251 226 52 324 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=46900 $D=1
M252 325 52 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=42270 $D=1
M253 326 52 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=46900 $D=1
M254 6 53 327 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=42270 $D=1
M255 7 53 328 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=46900 $D=1
M256 329 54 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=42270 $D=1
M257 330 54 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=46900 $D=1
M258 331 53 211 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=42270 $D=1
M259 332 53 212 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=46900 $D=1
M260 6 331 710 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=42270 $D=1
M261 7 332 711 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=46900 $D=1
M262 333 710 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=42270 $D=1
M263 334 711 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=46900 $D=1
M264 331 327 333 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=42270 $D=1
M265 332 328 334 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=46900 $D=1
M266 333 54 221 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=42270 $D=1
M267 334 54 222 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=46900 $D=1
M268 225 55 333 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=42270 $D=1
M269 226 55 334 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=46900 $D=1
M270 335 55 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=42270 $D=1
M271 336 55 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=46900 $D=1
M272 6 56 337 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=42270 $D=1
M273 7 56 338 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=46900 $D=1
M274 339 57 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=42270 $D=1
M275 340 57 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=46900 $D=1
M276 341 56 211 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=42270 $D=1
M277 342 56 212 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=46900 $D=1
M278 6 341 712 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=42270 $D=1
M279 7 342 713 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=46900 $D=1
M280 343 712 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=42270 $D=1
M281 344 713 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=46900 $D=1
M282 341 337 343 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=42270 $D=1
M283 342 338 344 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=46900 $D=1
M284 343 57 221 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=42270 $D=1
M285 344 57 222 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=46900 $D=1
M286 225 58 343 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=42270 $D=1
M287 226 58 344 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=46900 $D=1
M288 345 58 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=42270 $D=1
M289 346 58 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=46900 $D=1
M290 6 59 347 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=42270 $D=1
M291 7 59 348 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=46900 $D=1
M292 349 60 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=42270 $D=1
M293 350 60 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=46900 $D=1
M294 351 59 211 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=42270 $D=1
M295 352 59 212 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=46900 $D=1
M296 6 351 714 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=42270 $D=1
M297 7 352 715 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=46900 $D=1
M298 353 714 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=42270 $D=1
M299 354 715 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=46900 $D=1
M300 351 347 353 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=42270 $D=1
M301 352 348 354 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=46900 $D=1
M302 353 60 221 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=42270 $D=1
M303 354 60 222 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=46900 $D=1
M304 225 61 353 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=42270 $D=1
M305 226 61 354 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=46900 $D=1
M306 355 61 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=42270 $D=1
M307 356 61 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=46900 $D=1
M308 6 62 357 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=42270 $D=1
M309 7 62 358 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=46900 $D=1
M310 359 63 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=42270 $D=1
M311 360 63 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=46900 $D=1
M312 361 62 211 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=42270 $D=1
M313 362 62 212 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=46900 $D=1
M314 6 361 716 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=42270 $D=1
M315 7 362 717 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=46900 $D=1
M316 363 716 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=42270 $D=1
M317 364 717 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=46900 $D=1
M318 361 357 363 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=42270 $D=1
M319 362 358 364 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=46900 $D=1
M320 363 63 221 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=42270 $D=1
M321 364 63 222 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=46900 $D=1
M322 225 64 363 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=42270 $D=1
M323 226 64 364 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=46900 $D=1
M324 365 64 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=42270 $D=1
M325 366 64 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=46900 $D=1
M326 6 65 367 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=42270 $D=1
M327 7 65 368 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=46900 $D=1
M328 369 66 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=42270 $D=1
M329 370 66 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=46900 $D=1
M330 371 65 211 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=42270 $D=1
M331 372 65 212 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=46900 $D=1
M332 6 371 718 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=42270 $D=1
M333 7 372 719 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=46900 $D=1
M334 373 718 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=42270 $D=1
M335 374 719 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=46900 $D=1
M336 371 367 373 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=42270 $D=1
M337 372 368 374 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=46900 $D=1
M338 373 66 221 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=42270 $D=1
M339 374 66 222 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=46900 $D=1
M340 225 67 373 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=42270 $D=1
M341 226 67 374 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=46900 $D=1
M342 375 67 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=42270 $D=1
M343 376 67 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=46900 $D=1
M344 6 68 377 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=42270 $D=1
M345 7 68 378 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=46900 $D=1
M346 379 69 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=42270 $D=1
M347 380 69 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=46900 $D=1
M348 381 68 211 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=42270 $D=1
M349 382 68 212 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=46900 $D=1
M350 6 381 720 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=42270 $D=1
M351 7 382 721 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=46900 $D=1
M352 383 720 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=42270 $D=1
M353 384 721 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=46900 $D=1
M354 381 377 383 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=42270 $D=1
M355 382 378 384 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=46900 $D=1
M356 383 69 221 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=42270 $D=1
M357 384 69 222 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=46900 $D=1
M358 225 70 383 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=42270 $D=1
M359 226 70 384 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=46900 $D=1
M360 385 70 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=42270 $D=1
M361 386 70 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=46900 $D=1
M362 6 71 387 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=42270 $D=1
M363 7 71 388 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=46900 $D=1
M364 389 72 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=42270 $D=1
M365 390 72 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=46900 $D=1
M366 391 71 211 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=42270 $D=1
M367 392 71 212 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=46900 $D=1
M368 6 391 722 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=42270 $D=1
M369 7 392 723 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=46900 $D=1
M370 393 722 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=42270 $D=1
M371 394 723 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=46900 $D=1
M372 391 387 393 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=42270 $D=1
M373 392 388 394 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=46900 $D=1
M374 393 72 221 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=42270 $D=1
M375 394 72 222 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=46900 $D=1
M376 225 73 393 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=42270 $D=1
M377 226 73 394 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=46900 $D=1
M378 395 73 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=42270 $D=1
M379 396 73 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=46900 $D=1
M380 6 74 397 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=42270 $D=1
M381 7 74 398 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=46900 $D=1
M382 399 75 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=42270 $D=1
M383 400 75 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=46900 $D=1
M384 401 74 211 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=42270 $D=1
M385 402 74 212 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=46900 $D=1
M386 6 401 724 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=42270 $D=1
M387 7 402 725 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=46900 $D=1
M388 403 724 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=42270 $D=1
M389 404 725 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=46900 $D=1
M390 401 397 403 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=42270 $D=1
M391 402 398 404 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=46900 $D=1
M392 403 75 221 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=42270 $D=1
M393 404 75 222 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=46900 $D=1
M394 225 76 403 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=42270 $D=1
M395 226 76 404 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=46900 $D=1
M396 405 76 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=42270 $D=1
M397 406 76 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=46900 $D=1
M398 6 77 407 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=42270 $D=1
M399 7 77 408 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=46900 $D=1
M400 409 78 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=42270 $D=1
M401 410 78 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=46900 $D=1
M402 411 77 211 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=42270 $D=1
M403 412 77 212 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=46900 $D=1
M404 6 411 726 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=42270 $D=1
M405 7 412 727 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=46900 $D=1
M406 413 726 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=42270 $D=1
M407 414 727 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=46900 $D=1
M408 411 407 413 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=42270 $D=1
M409 412 408 414 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=46900 $D=1
M410 413 78 221 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=42270 $D=1
M411 414 78 222 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=46900 $D=1
M412 225 79 413 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=42270 $D=1
M413 226 79 414 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=46900 $D=1
M414 415 79 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=42270 $D=1
M415 416 79 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=46900 $D=1
M416 6 80 417 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=42270 $D=1
M417 7 80 418 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=46900 $D=1
M418 419 81 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=42270 $D=1
M419 420 81 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=46900 $D=1
M420 421 80 211 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=42270 $D=1
M421 422 80 212 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=46900 $D=1
M422 6 421 728 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=42270 $D=1
M423 7 422 729 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=46900 $D=1
M424 423 728 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=42270 $D=1
M425 424 729 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=46900 $D=1
M426 421 417 423 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=42270 $D=1
M427 422 418 424 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=46900 $D=1
M428 423 81 221 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=42270 $D=1
M429 424 81 222 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=46900 $D=1
M430 225 82 423 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=42270 $D=1
M431 226 82 424 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=46900 $D=1
M432 425 82 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=42270 $D=1
M433 426 82 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=46900 $D=1
M434 6 83 427 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=42270 $D=1
M435 7 83 428 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=46900 $D=1
M436 429 84 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=42270 $D=1
M437 430 84 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=46900 $D=1
M438 431 83 211 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=42270 $D=1
M439 432 83 212 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=46900 $D=1
M440 6 431 730 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=42270 $D=1
M441 7 432 731 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=46900 $D=1
M442 433 730 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=42270 $D=1
M443 434 731 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=46900 $D=1
M444 431 427 433 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=42270 $D=1
M445 432 428 434 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=46900 $D=1
M446 433 84 221 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=42270 $D=1
M447 434 84 222 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=46900 $D=1
M448 225 85 433 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=42270 $D=1
M449 226 85 434 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=46900 $D=1
M450 435 85 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=42270 $D=1
M451 436 85 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=46900 $D=1
M452 6 86 437 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=42270 $D=1
M453 7 86 438 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=46900 $D=1
M454 439 87 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=42270 $D=1
M455 440 87 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=46900 $D=1
M456 441 86 211 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=42270 $D=1
M457 442 86 212 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=46900 $D=1
M458 6 441 732 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=42270 $D=1
M459 7 442 733 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=46900 $D=1
M460 443 732 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=42270 $D=1
M461 444 733 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=46900 $D=1
M462 441 437 443 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=42270 $D=1
M463 442 438 444 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=46900 $D=1
M464 443 87 221 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=42270 $D=1
M465 444 87 222 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=46900 $D=1
M466 225 88 443 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=42270 $D=1
M467 226 88 444 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=46900 $D=1
M468 445 88 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=42270 $D=1
M469 446 88 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=46900 $D=1
M470 6 89 447 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=42270 $D=1
M471 7 89 448 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=46900 $D=1
M472 449 90 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=42270 $D=1
M473 450 90 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=46900 $D=1
M474 451 89 211 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=42270 $D=1
M475 452 89 212 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=46900 $D=1
M476 6 451 734 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=42270 $D=1
M477 7 452 735 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=46900 $D=1
M478 453 734 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=42270 $D=1
M479 454 735 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=46900 $D=1
M480 451 447 453 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=42270 $D=1
M481 452 448 454 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=46900 $D=1
M482 453 90 221 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=42270 $D=1
M483 454 90 222 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=46900 $D=1
M484 225 91 453 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=42270 $D=1
M485 226 91 454 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=46900 $D=1
M486 455 91 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=42270 $D=1
M487 456 91 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=46900 $D=1
M488 6 92 457 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=42270 $D=1
M489 7 92 458 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=46900 $D=1
M490 459 93 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=42270 $D=1
M491 460 93 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=46900 $D=1
M492 461 92 211 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=42270 $D=1
M493 462 92 212 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=46900 $D=1
M494 6 461 736 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=42270 $D=1
M495 7 462 737 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=46900 $D=1
M496 463 736 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=42270 $D=1
M497 464 737 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=46900 $D=1
M498 461 457 463 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=42270 $D=1
M499 462 458 464 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=46900 $D=1
M500 463 93 221 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=42270 $D=1
M501 464 93 222 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=46900 $D=1
M502 225 94 463 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=42270 $D=1
M503 226 94 464 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=46900 $D=1
M504 465 94 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=42270 $D=1
M505 466 94 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=46900 $D=1
M506 6 95 467 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=42270 $D=1
M507 7 95 468 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=46900 $D=1
M508 469 96 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=42270 $D=1
M509 470 96 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=46900 $D=1
M510 471 95 211 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=42270 $D=1
M511 472 95 212 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=46900 $D=1
M512 6 471 738 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=42270 $D=1
M513 7 472 739 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=46900 $D=1
M514 473 738 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=42270 $D=1
M515 474 739 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=46900 $D=1
M516 471 467 473 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=42270 $D=1
M517 472 468 474 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=46900 $D=1
M518 473 96 221 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=42270 $D=1
M519 474 96 222 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=46900 $D=1
M520 225 97 473 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=42270 $D=1
M521 226 97 474 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=46900 $D=1
M522 475 97 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=42270 $D=1
M523 476 97 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=46900 $D=1
M524 6 98 477 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=42270 $D=1
M525 7 98 478 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=46900 $D=1
M526 479 99 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=42270 $D=1
M527 480 99 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=46900 $D=1
M528 481 98 211 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=42270 $D=1
M529 482 98 212 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=46900 $D=1
M530 6 481 740 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=42270 $D=1
M531 7 482 741 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=46900 $D=1
M532 483 740 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=42270 $D=1
M533 484 741 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=46900 $D=1
M534 481 477 483 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=42270 $D=1
M535 482 478 484 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=46900 $D=1
M536 483 99 221 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=42270 $D=1
M537 484 99 222 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=46900 $D=1
M538 225 100 483 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=42270 $D=1
M539 226 100 484 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=46900 $D=1
M540 485 100 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=42270 $D=1
M541 486 100 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=46900 $D=1
M542 6 101 487 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=42270 $D=1
M543 7 101 488 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=46900 $D=1
M544 489 102 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=42270 $D=1
M545 490 102 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=46900 $D=1
M546 491 101 211 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=42270 $D=1
M547 492 101 212 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=46900 $D=1
M548 6 491 742 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=42270 $D=1
M549 7 492 743 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=46900 $D=1
M550 493 742 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=42270 $D=1
M551 494 743 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=46900 $D=1
M552 491 487 493 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=42270 $D=1
M553 492 488 494 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=46900 $D=1
M554 493 102 221 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=42270 $D=1
M555 494 102 222 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=46900 $D=1
M556 225 103 493 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=42270 $D=1
M557 226 103 494 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=46900 $D=1
M558 495 103 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=42270 $D=1
M559 496 103 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=46900 $D=1
M560 6 104 497 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=42270 $D=1
M561 7 104 498 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=46900 $D=1
M562 499 105 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=42270 $D=1
M563 500 105 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=46900 $D=1
M564 501 104 211 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=42270 $D=1
M565 502 104 212 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=46900 $D=1
M566 6 501 744 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=42270 $D=1
M567 7 502 745 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=46900 $D=1
M568 503 744 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=42270 $D=1
M569 504 745 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=46900 $D=1
M570 501 497 503 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=42270 $D=1
M571 502 498 504 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=46900 $D=1
M572 503 105 221 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=42270 $D=1
M573 504 105 222 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=46900 $D=1
M574 225 106 503 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=42270 $D=1
M575 226 106 504 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=46900 $D=1
M576 505 106 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=42270 $D=1
M577 506 106 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=46900 $D=1
M578 6 107 507 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=42270 $D=1
M579 7 107 508 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=46900 $D=1
M580 509 108 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=42270 $D=1
M581 510 108 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=46900 $D=1
M582 511 107 211 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=42270 $D=1
M583 512 107 212 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=46900 $D=1
M584 6 511 746 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=42270 $D=1
M585 7 512 747 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=46900 $D=1
M586 513 746 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=42270 $D=1
M587 514 747 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=46900 $D=1
M588 511 507 513 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=42270 $D=1
M589 512 508 514 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=46900 $D=1
M590 513 108 221 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=42270 $D=1
M591 514 108 222 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=46900 $D=1
M592 225 109 513 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=42270 $D=1
M593 226 109 514 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=46900 $D=1
M594 515 109 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=42270 $D=1
M595 516 109 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=46900 $D=1
M596 6 110 517 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=42270 $D=1
M597 7 110 518 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=46900 $D=1
M598 519 111 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=42270 $D=1
M599 520 111 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=46900 $D=1
M600 521 110 211 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=42270 $D=1
M601 522 110 212 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=46900 $D=1
M602 6 521 748 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=42270 $D=1
M603 7 522 749 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=46900 $D=1
M604 523 748 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=42270 $D=1
M605 524 749 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=46900 $D=1
M606 521 517 523 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=42270 $D=1
M607 522 518 524 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=46900 $D=1
M608 523 111 221 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=42270 $D=1
M609 524 111 222 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=46900 $D=1
M610 225 112 523 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=42270 $D=1
M611 226 112 524 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=46900 $D=1
M612 525 112 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=42270 $D=1
M613 526 112 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=46900 $D=1
M614 6 113 527 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=42270 $D=1
M615 7 113 528 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=46900 $D=1
M616 529 114 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=42270 $D=1
M617 530 114 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=46900 $D=1
M618 6 114 221 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=42270 $D=1
M619 7 114 222 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=46900 $D=1
M620 225 113 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=42270 $D=1
M621 226 113 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=46900 $D=1
M622 6 533 531 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=42270 $D=1
M623 7 534 532 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=46900 $D=1
M624 533 115 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=42270 $D=1
M625 534 115 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=46900 $D=1
M626 750 221 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=42270 $D=1
M627 751 222 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=46900 $D=1
M628 535 531 750 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=42270 $D=1
M629 536 532 751 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=46900 $D=1
M630 6 535 537 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=42270 $D=1
M631 7 536 538 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=46900 $D=1
M632 752 537 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=42270 $D=1
M633 753 538 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=46900 $D=1
M634 535 533 752 6 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=42270 $D=1
M635 536 534 753 7 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=46900 $D=1
M636 6 541 539 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=42270 $D=1
M637 7 542 540 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=46900 $D=1
M638 541 115 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=42270 $D=1
M639 542 115 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=46900 $D=1
M640 754 225 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=42270 $D=1
M641 755 226 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=46900 $D=1
M642 543 539 754 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=42270 $D=1
M643 544 540 755 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=46900 $D=1
M644 6 543 116 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=42270 $D=1
M645 7 544 117 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=46900 $D=1
M646 756 116 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=42270 $D=1
M647 757 117 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=46900 $D=1
M648 543 541 756 6 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=42270 $D=1
M649 544 542 757 7 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=46900 $D=1
M650 545 118 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=42270 $D=1
M651 546 118 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=46900 $D=1
M652 547 545 537 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=42270 $D=1
M653 548 546 538 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=46900 $D=1
M654 119 118 547 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=42270 $D=1
M655 120 118 548 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=46900 $D=1
M656 549 121 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=42270 $D=1
M657 550 121 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=46900 $D=1
M658 551 549 116 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=42270 $D=1
M659 552 550 117 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=46900 $D=1
M660 758 121 551 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=42270 $D=1
M661 759 121 552 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=46900 $D=1
M662 6 116 758 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=42270 $D=1
M663 7 117 759 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=46900 $D=1
M664 553 122 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=42270 $D=1
M665 554 122 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=46900 $D=1
M666 555 553 551 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=42270 $D=1
M667 556 554 552 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=46900 $D=1
M668 12 122 555 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=42270 $D=1
M669 13 122 556 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=46900 $D=1
M670 559 557 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=42270 $D=1
M671 560 558 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=46900 $D=1
M672 6 563 561 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=42270 $D=1
M673 7 564 562 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=46900 $D=1
M674 565 547 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=42270 $D=1
M675 566 548 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=46900 $D=1
M676 563 565 557 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=42270 $D=1
M677 564 566 558 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=46900 $D=1
M678 559 547 563 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=42270 $D=1
M679 560 548 564 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=46900 $D=1
M680 567 561 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=42270 $D=1
M681 568 562 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=46900 $D=1
M682 123 567 555 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=42270 $D=1
M683 557 568 556 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=46900 $D=1
M684 547 561 123 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=42270 $D=1
M685 548 562 557 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=46900 $D=1
M686 569 123 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=42270 $D=1
M687 570 557 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=46900 $D=1
M688 571 561 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=42270 $D=1
M689 572 562 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=46900 $D=1
M690 573 571 569 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=42270 $D=1
M691 574 572 570 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=46900 $D=1
M692 555 561 573 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=42270 $D=1
M693 556 562 574 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=46900 $D=1
M694 575 547 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=42270 $D=1
M695 576 548 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=46900 $D=1
M696 6 555 575 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=42270 $D=1
M697 7 556 576 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=46900 $D=1
M698 577 573 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=42270 $D=1
M699 578 574 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=46900 $D=1
M700 786 547 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=42270 $D=1
M701 787 548 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=46900 $D=1
M702 579 555 786 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=42270 $D=1
M703 580 556 787 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=46900 $D=1
M704 788 547 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=42270 $D=1
M705 789 548 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=46900 $D=1
M706 581 555 788 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=42270 $D=1
M707 582 556 789 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=46900 $D=1
M708 585 547 583 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=42270 $D=1
M709 586 548 584 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=46900 $D=1
M710 583 555 585 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=42270 $D=1
M711 584 556 586 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=46900 $D=1
M712 6 581 583 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=42270 $D=1
M713 7 582 584 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=46900 $D=1
M714 587 128 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=42270 $D=1
M715 588 128 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=46900 $D=1
M716 589 587 575 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=42270 $D=1
M717 590 588 576 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=46900 $D=1
M718 579 128 589 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=42270 $D=1
M719 580 128 590 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=46900 $D=1
M720 591 587 577 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=42270 $D=1
M721 592 588 578 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=46900 $D=1
M722 585 128 591 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=42270 $D=1
M723 586 128 592 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=46900 $D=1
M724 593 129 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=42270 $D=1
M725 594 129 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=46900 $D=1
M726 595 593 591 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=42270 $D=1
M727 596 594 592 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=46900 $D=1
M728 589 129 595 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=42270 $D=1
M729 590 129 596 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=46900 $D=1
M730 14 595 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=42270 $D=1
M731 15 596 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=46900 $D=1
M732 597 130 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=42270 $D=1
M733 598 130 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=46900 $D=1
M734 599 597 131 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=42270 $D=1
M735 600 598 132 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=46900 $D=1
M736 133 130 599 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=42270 $D=1
M737 134 130 600 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=46900 $D=1
M738 601 130 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=42270 $D=1
M739 602 130 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=46900 $D=1
M740 604 601 135 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=42270 $D=1
M741 605 602 137 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=46900 $D=1
M742 138 130 604 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=42270 $D=1
M743 136 130 605 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=46900 $D=1
M744 606 130 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=42270 $D=1
M745 607 130 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=46900 $D=1
M746 608 606 127 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=42270 $D=1
M747 609 607 126 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=46900 $D=1
M748 139 130 608 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=42270 $D=1
M749 140 130 609 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=46900 $D=1
M750 610 130 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=42270 $D=1
M751 611 130 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=46900 $D=1
M752 612 610 141 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=42270 $D=1
M753 613 611 142 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=46900 $D=1
M754 143 130 612 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=42270 $D=1
M755 144 130 613 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=46900 $D=1
M756 614 130 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=42270 $D=1
M757 615 130 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=46900 $D=1
M758 616 614 145 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=42270 $D=1
M759 617 615 146 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=46900 $D=1
M760 147 130 616 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=42270 $D=1
M761 147 130 617 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=46900 $D=1
M762 6 547 768 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=42270 $D=1
M763 7 548 769 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=46900 $D=1
M764 134 768 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=42270 $D=1
M765 131 769 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=46900 $D=1
M766 618 148 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=42270 $D=1
M767 619 148 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=46900 $D=1
M768 149 618 134 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=42270 $D=1
M769 150 619 131 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=46900 $D=1
M770 599 148 149 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=42270 $D=1
M771 600 148 150 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=46900 $D=1
M772 620 151 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=42270 $D=1
M773 621 151 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=46900 $D=1
M774 152 620 149 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=42270 $D=1
M775 125 621 150 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=46900 $D=1
M776 604 151 152 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=42270 $D=1
M777 605 151 125 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=46900 $D=1
M778 622 153 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=42270 $D=1
M779 623 153 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=46900 $D=1
M780 154 622 152 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=42270 $D=1
M781 155 623 125 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=46900 $D=1
M782 608 153 154 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=42270 $D=1
M783 609 153 155 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=46900 $D=1
M784 624 156 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=42270 $D=1
M785 625 156 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=46900 $D=1
M786 157 624 154 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=42270 $D=1
M787 158 625 155 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=46900 $D=1
M788 612 156 157 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=42270 $D=1
M789 613 156 158 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=46900 $D=1
M790 626 159 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=42270 $D=1
M791 627 159 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=46900 $D=1
M792 16 626 157 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=42270 $D=1
M793 17 627 158 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=46900 $D=1
M794 616 159 16 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=42270 $D=1
M795 617 159 17 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=46900 $D=1
M796 628 160 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=42270 $D=1
M797 629 160 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=46900 $D=1
M798 630 628 116 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=42270 $D=1
M799 631 629 117 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=46900 $D=1
M800 12 160 630 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=42270 $D=1
M801 13 160 631 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=46900 $D=1
M802 790 537 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=42270 $D=1
M803 791 538 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=46900 $D=1
M804 632 630 790 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=42270 $D=1
M805 633 631 791 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=46900 $D=1
M806 636 537 634 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=42270 $D=1
M807 637 538 635 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=46900 $D=1
M808 634 630 636 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=42270 $D=1
M809 635 631 637 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=46900 $D=1
M810 6 632 634 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=42270 $D=1
M811 7 633 635 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=46900 $D=1
M812 792 161 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=42270 $D=1
M813 793 638 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=46900 $D=1
M814 770 636 792 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=42270 $D=1
M815 771 637 793 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=46900 $D=1
M816 638 770 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=42270 $D=1
M817 639 771 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=46900 $D=1
M818 640 537 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=42270 $D=1
M819 641 538 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=46900 $D=1
M820 6 642 640 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=42270 $D=1
M821 7 643 641 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=46900 $D=1
M822 642 630 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=42270 $D=1
M823 643 631 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=46900 $D=1
M824 794 640 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=42270 $D=1
M825 795 641 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=46900 $D=1
M826 644 161 794 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=42270 $D=1
M827 645 638 795 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=46900 $D=1
M828 647 162 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=42270 $D=1
M829 648 646 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=46900 $D=1
M830 796 644 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=42270 $D=1
M831 797 645 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=46900 $D=1
M832 646 647 796 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=42270 $D=1
M833 163 648 797 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=46900 $D=1
M834 650 649 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=42270 $D=1
M835 651 164 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=46900 $D=1
M836 6 654 652 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=42270 $D=1
M837 7 655 653 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=46900 $D=1
M838 656 119 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=42270 $D=1
M839 657 120 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=46900 $D=1
M840 654 656 649 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=42270 $D=1
M841 655 657 164 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=46900 $D=1
M842 650 119 654 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=42270 $D=1
M843 651 120 655 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=46900 $D=1
M844 658 652 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=42270 $D=1
M845 659 653 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=46900 $D=1
M846 165 658 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=42270 $D=1
M847 649 659 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=46900 $D=1
M848 119 652 165 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=42270 $D=1
M849 120 653 649 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=46900 $D=1
M850 660 165 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=42270 $D=1
M851 661 649 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=46900 $D=1
M852 662 652 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=42270 $D=1
M853 663 653 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=46900 $D=1
M854 199 662 660 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=42270 $D=1
M855 200 663 661 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=46900 $D=1
M856 6 652 199 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=42270 $D=1
M857 7 653 200 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=46900 $D=1
M858 664 166 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=42270 $D=1
M859 665 166 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=46900 $D=1
M860 666 664 199 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=42270 $D=1
M861 667 665 200 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=46900 $D=1
M862 14 166 666 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=42270 $D=1
M863 15 166 667 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=46900 $D=1
M864 668 167 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=42270 $D=1
M865 669 167 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=46900 $D=1
M866 167 668 666 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=42270 $D=1
M867 167 669 667 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=46900 $D=1
M868 6 167 167 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=42270 $D=1
M869 7 167 167 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=46900 $D=1
M870 670 115 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=42270 $D=1
M871 671 115 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=46900 $D=1
M872 6 670 672 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=42270 $D=1
M873 7 671 673 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=46900 $D=1
M874 674 115 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=42270 $D=1
M875 675 115 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=46900 $D=1
M876 676 670 167 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=42270 $D=1
M877 677 671 167 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=46900 $D=1
M878 6 676 772 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=42270 $D=1
M879 7 677 773 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=46900 $D=1
M880 678 772 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=42270 $D=1
M881 679 773 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=46900 $D=1
M882 676 672 678 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=42270 $D=1
M883 677 673 679 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=46900 $D=1
M884 680 115 678 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=42270 $D=1
M885 681 115 679 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=46900 $D=1
M886 6 684 682 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=42270 $D=1
M887 7 685 683 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=46900 $D=1
M888 684 115 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=42270 $D=1
M889 685 115 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=46900 $D=1
M890 774 680 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=42270 $D=1
M891 775 681 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=46900 $D=1
M892 686 682 774 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=42270 $D=1
M893 687 683 775 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=46900 $D=1
M894 6 686 119 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=42270 $D=1
M895 7 687 120 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=46900 $D=1
M896 776 119 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=42270 $D=1
M897 777 120 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=46900 $D=1
M898 686 684 776 6 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=42270 $D=1
M899 687 685 777 7 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=46900 $D=1
M900 175 1 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=43520 $D=0
M901 176 1 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=48150 $D=0
M902 177 1 2 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=43520 $D=0
M903 178 1 3 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=48150 $D=0
M904 6 175 177 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=43520 $D=0
M905 7 176 178 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=48150 $D=0
M906 179 1 4 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=43520 $D=0
M907 180 1 4 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=48150 $D=0
M908 5 175 179 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=43520 $D=0
M909 5 176 180 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=48150 $D=0
M910 181 1 6 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=43520 $D=0
M911 182 1 7 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=48150 $D=0
M912 6 175 181 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=43520 $D=0
M913 7 176 182 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=48150 $D=0
M914 185 9 181 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=43520 $D=0
M915 186 9 182 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=48150 $D=0
M916 183 9 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=43520 $D=0
M917 184 9 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=48150 $D=0
M918 187 9 179 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=43520 $D=0
M919 188 9 180 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=48150 $D=0
M920 177 183 187 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=43520 $D=0
M921 178 184 188 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=48150 $D=0
M922 189 10 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=43520 $D=0
M923 190 10 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=48150 $D=0
M924 191 10 187 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=43520 $D=0
M925 192 10 188 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=48150 $D=0
M926 185 189 191 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=43520 $D=0
M927 186 190 192 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=48150 $D=0
M928 193 11 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=43520 $D=0
M929 194 11 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=48150 $D=0
M930 195 11 6 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=43520 $D=0
M931 196 11 7 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=48150 $D=0
M932 12 193 195 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=43520 $D=0
M933 13 194 196 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=48150 $D=0
M934 197 11 14 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=43520 $D=0
M935 198 11 15 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=48150 $D=0
M936 16 193 197 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=43520 $D=0
M937 17 194 198 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=48150 $D=0
M938 201 11 199 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=43520 $D=0
M939 202 11 200 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=48150 $D=0
M940 191 193 201 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=43520 $D=0
M941 192 194 202 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=48150 $D=0
M942 205 18 201 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=43520 $D=0
M943 206 18 202 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=48150 $D=0
M944 203 18 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=43520 $D=0
M945 204 18 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=48150 $D=0
M946 207 18 197 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=43520 $D=0
M947 208 18 198 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=48150 $D=0
M948 195 203 207 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=43520 $D=0
M949 196 204 208 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=48150 $D=0
M950 209 19 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=43520 $D=0
M951 210 19 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=48150 $D=0
M952 211 19 207 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=43520 $D=0
M953 212 19 208 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=48150 $D=0
M954 205 209 211 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=43520 $D=0
M955 206 210 212 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=48150 $D=0
M956 168 20 213 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=43520 $D=0
M957 169 20 214 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=48150 $D=0
M958 215 21 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=43520 $D=0
M959 216 21 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=48150 $D=0
M960 217 213 211 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=43520 $D=0
M961 218 214 212 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=48150 $D=0
M962 168 217 688 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=43520 $D=0
M963 169 218 689 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=48150 $D=0
M964 219 688 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=43520 $D=0
M965 220 689 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=48150 $D=0
M966 217 20 219 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=43520 $D=0
M967 218 20 220 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=48150 $D=0
M968 219 215 221 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=43520 $D=0
M969 220 216 222 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=48150 $D=0
M970 225 223 219 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=43520 $D=0
M971 226 224 220 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=48150 $D=0
M972 223 22 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=43520 $D=0
M973 224 22 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=48150 $D=0
M974 168 23 227 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=43520 $D=0
M975 169 23 228 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=48150 $D=0
M976 229 24 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=43520 $D=0
M977 230 24 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=48150 $D=0
M978 231 227 211 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=43520 $D=0
M979 232 228 212 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=48150 $D=0
M980 168 231 690 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=43520 $D=0
M981 169 232 691 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=48150 $D=0
M982 233 690 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=43520 $D=0
M983 234 691 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=48150 $D=0
M984 231 23 233 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=43520 $D=0
M985 232 23 234 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=48150 $D=0
M986 233 229 221 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=43520 $D=0
M987 234 230 222 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=48150 $D=0
M988 225 235 233 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=43520 $D=0
M989 226 236 234 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=48150 $D=0
M990 235 25 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=43520 $D=0
M991 236 25 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=48150 $D=0
M992 168 26 237 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=43520 $D=0
M993 169 26 238 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=48150 $D=0
M994 239 27 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=43520 $D=0
M995 240 27 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=48150 $D=0
M996 241 237 211 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=43520 $D=0
M997 242 238 212 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=48150 $D=0
M998 168 241 692 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=43520 $D=0
M999 169 242 693 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=48150 $D=0
M1000 243 692 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=43520 $D=0
M1001 244 693 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=48150 $D=0
M1002 241 26 243 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=43520 $D=0
M1003 242 26 244 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=48150 $D=0
M1004 243 239 221 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=43520 $D=0
M1005 244 240 222 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=48150 $D=0
M1006 225 245 243 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=43520 $D=0
M1007 226 246 244 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=48150 $D=0
M1008 245 28 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=43520 $D=0
M1009 246 28 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=48150 $D=0
M1010 168 29 247 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=43520 $D=0
M1011 169 29 248 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=48150 $D=0
M1012 249 30 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=43520 $D=0
M1013 250 30 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=48150 $D=0
M1014 251 247 211 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=43520 $D=0
M1015 252 248 212 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=48150 $D=0
M1016 168 251 694 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=43520 $D=0
M1017 169 252 695 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=48150 $D=0
M1018 253 694 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=43520 $D=0
M1019 254 695 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=48150 $D=0
M1020 251 29 253 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=43520 $D=0
M1021 252 29 254 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=48150 $D=0
M1022 253 249 221 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=43520 $D=0
M1023 254 250 222 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=48150 $D=0
M1024 225 255 253 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=43520 $D=0
M1025 226 256 254 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=48150 $D=0
M1026 255 31 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=43520 $D=0
M1027 256 31 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=48150 $D=0
M1028 168 32 257 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=43520 $D=0
M1029 169 32 258 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=48150 $D=0
M1030 259 33 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=43520 $D=0
M1031 260 33 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=48150 $D=0
M1032 261 257 211 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=43520 $D=0
M1033 262 258 212 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=48150 $D=0
M1034 168 261 696 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=43520 $D=0
M1035 169 262 697 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=48150 $D=0
M1036 263 696 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=43520 $D=0
M1037 264 697 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=48150 $D=0
M1038 261 32 263 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=43520 $D=0
M1039 262 32 264 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=48150 $D=0
M1040 263 259 221 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=43520 $D=0
M1041 264 260 222 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=48150 $D=0
M1042 225 265 263 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=43520 $D=0
M1043 226 266 264 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=48150 $D=0
M1044 265 34 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=43520 $D=0
M1045 266 34 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=48150 $D=0
M1046 168 35 267 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=43520 $D=0
M1047 169 35 268 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=48150 $D=0
M1048 269 36 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=43520 $D=0
M1049 270 36 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=48150 $D=0
M1050 271 267 211 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=43520 $D=0
M1051 272 268 212 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=48150 $D=0
M1052 168 271 698 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=43520 $D=0
M1053 169 272 699 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=48150 $D=0
M1054 273 698 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=43520 $D=0
M1055 274 699 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=48150 $D=0
M1056 271 35 273 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=43520 $D=0
M1057 272 35 274 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=48150 $D=0
M1058 273 269 221 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=43520 $D=0
M1059 274 270 222 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=48150 $D=0
M1060 225 275 273 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=43520 $D=0
M1061 226 276 274 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=48150 $D=0
M1062 275 37 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=43520 $D=0
M1063 276 37 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=48150 $D=0
M1064 168 38 277 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=43520 $D=0
M1065 169 38 278 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=48150 $D=0
M1066 279 39 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=43520 $D=0
M1067 280 39 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=48150 $D=0
M1068 281 277 211 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=43520 $D=0
M1069 282 278 212 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=48150 $D=0
M1070 168 281 700 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=43520 $D=0
M1071 169 282 701 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=48150 $D=0
M1072 283 700 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=43520 $D=0
M1073 284 701 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=48150 $D=0
M1074 281 38 283 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=43520 $D=0
M1075 282 38 284 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=48150 $D=0
M1076 283 279 221 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=43520 $D=0
M1077 284 280 222 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=48150 $D=0
M1078 225 285 283 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=43520 $D=0
M1079 226 286 284 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=48150 $D=0
M1080 285 40 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=43520 $D=0
M1081 286 40 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=48150 $D=0
M1082 168 41 287 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=43520 $D=0
M1083 169 41 288 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=48150 $D=0
M1084 289 42 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=43520 $D=0
M1085 290 42 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=48150 $D=0
M1086 291 287 211 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=43520 $D=0
M1087 292 288 212 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=48150 $D=0
M1088 168 291 702 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=43520 $D=0
M1089 169 292 703 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=48150 $D=0
M1090 293 702 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=43520 $D=0
M1091 294 703 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=48150 $D=0
M1092 291 41 293 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=43520 $D=0
M1093 292 41 294 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=48150 $D=0
M1094 293 289 221 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=43520 $D=0
M1095 294 290 222 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=48150 $D=0
M1096 225 295 293 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=43520 $D=0
M1097 226 296 294 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=48150 $D=0
M1098 295 43 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=43520 $D=0
M1099 296 43 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=48150 $D=0
M1100 168 44 297 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=43520 $D=0
M1101 169 44 298 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=48150 $D=0
M1102 299 45 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=43520 $D=0
M1103 300 45 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=48150 $D=0
M1104 301 297 211 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=43520 $D=0
M1105 302 298 212 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=48150 $D=0
M1106 168 301 704 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=43520 $D=0
M1107 169 302 705 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=48150 $D=0
M1108 303 704 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=43520 $D=0
M1109 304 705 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=48150 $D=0
M1110 301 44 303 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=43520 $D=0
M1111 302 44 304 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=48150 $D=0
M1112 303 299 221 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=43520 $D=0
M1113 304 300 222 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=48150 $D=0
M1114 225 305 303 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=43520 $D=0
M1115 226 306 304 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=48150 $D=0
M1116 305 46 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=43520 $D=0
M1117 306 46 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=48150 $D=0
M1118 168 47 307 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=43520 $D=0
M1119 169 47 308 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=48150 $D=0
M1120 309 48 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=43520 $D=0
M1121 310 48 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=48150 $D=0
M1122 311 307 211 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=43520 $D=0
M1123 312 308 212 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=48150 $D=0
M1124 168 311 706 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=43520 $D=0
M1125 169 312 707 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=48150 $D=0
M1126 313 706 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=43520 $D=0
M1127 314 707 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=48150 $D=0
M1128 311 47 313 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=43520 $D=0
M1129 312 47 314 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=48150 $D=0
M1130 313 309 221 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=43520 $D=0
M1131 314 310 222 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=48150 $D=0
M1132 225 315 313 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=43520 $D=0
M1133 226 316 314 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=48150 $D=0
M1134 315 49 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=43520 $D=0
M1135 316 49 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=48150 $D=0
M1136 168 50 317 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=43520 $D=0
M1137 169 50 318 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=48150 $D=0
M1138 319 51 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=43520 $D=0
M1139 320 51 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=48150 $D=0
M1140 321 317 211 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=43520 $D=0
M1141 322 318 212 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=48150 $D=0
M1142 168 321 708 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=43520 $D=0
M1143 169 322 709 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=48150 $D=0
M1144 323 708 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=43520 $D=0
M1145 324 709 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=48150 $D=0
M1146 321 50 323 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=43520 $D=0
M1147 322 50 324 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=48150 $D=0
M1148 323 319 221 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=43520 $D=0
M1149 324 320 222 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=48150 $D=0
M1150 225 325 323 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=43520 $D=0
M1151 226 326 324 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=48150 $D=0
M1152 325 52 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=43520 $D=0
M1153 326 52 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=48150 $D=0
M1154 168 53 327 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=43520 $D=0
M1155 169 53 328 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=48150 $D=0
M1156 329 54 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=43520 $D=0
M1157 330 54 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=48150 $D=0
M1158 331 327 211 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=43520 $D=0
M1159 332 328 212 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=48150 $D=0
M1160 168 331 710 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=43520 $D=0
M1161 169 332 711 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=48150 $D=0
M1162 333 710 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=43520 $D=0
M1163 334 711 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=48150 $D=0
M1164 331 53 333 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=43520 $D=0
M1165 332 53 334 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=48150 $D=0
M1166 333 329 221 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=43520 $D=0
M1167 334 330 222 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=48150 $D=0
M1168 225 335 333 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=43520 $D=0
M1169 226 336 334 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=48150 $D=0
M1170 335 55 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=43520 $D=0
M1171 336 55 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=48150 $D=0
M1172 168 56 337 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=43520 $D=0
M1173 169 56 338 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=48150 $D=0
M1174 339 57 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=43520 $D=0
M1175 340 57 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=48150 $D=0
M1176 341 337 211 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=43520 $D=0
M1177 342 338 212 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=48150 $D=0
M1178 168 341 712 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=43520 $D=0
M1179 169 342 713 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=48150 $D=0
M1180 343 712 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=43520 $D=0
M1181 344 713 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=48150 $D=0
M1182 341 56 343 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=43520 $D=0
M1183 342 56 344 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=48150 $D=0
M1184 343 339 221 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=43520 $D=0
M1185 344 340 222 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=48150 $D=0
M1186 225 345 343 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=43520 $D=0
M1187 226 346 344 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=48150 $D=0
M1188 345 58 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=43520 $D=0
M1189 346 58 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=48150 $D=0
M1190 168 59 347 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=43520 $D=0
M1191 169 59 348 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=48150 $D=0
M1192 349 60 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=43520 $D=0
M1193 350 60 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=48150 $D=0
M1194 351 347 211 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=43520 $D=0
M1195 352 348 212 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=48150 $D=0
M1196 168 351 714 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=43520 $D=0
M1197 169 352 715 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=48150 $D=0
M1198 353 714 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=43520 $D=0
M1199 354 715 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=48150 $D=0
M1200 351 59 353 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=43520 $D=0
M1201 352 59 354 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=48150 $D=0
M1202 353 349 221 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=43520 $D=0
M1203 354 350 222 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=48150 $D=0
M1204 225 355 353 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=43520 $D=0
M1205 226 356 354 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=48150 $D=0
M1206 355 61 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=43520 $D=0
M1207 356 61 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=48150 $D=0
M1208 168 62 357 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=43520 $D=0
M1209 169 62 358 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=48150 $D=0
M1210 359 63 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=43520 $D=0
M1211 360 63 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=48150 $D=0
M1212 361 357 211 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=43520 $D=0
M1213 362 358 212 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=48150 $D=0
M1214 168 361 716 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=43520 $D=0
M1215 169 362 717 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=48150 $D=0
M1216 363 716 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=43520 $D=0
M1217 364 717 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=48150 $D=0
M1218 361 62 363 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=43520 $D=0
M1219 362 62 364 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=48150 $D=0
M1220 363 359 221 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=43520 $D=0
M1221 364 360 222 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=48150 $D=0
M1222 225 365 363 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=43520 $D=0
M1223 226 366 364 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=48150 $D=0
M1224 365 64 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=43520 $D=0
M1225 366 64 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=48150 $D=0
M1226 168 65 367 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=43520 $D=0
M1227 169 65 368 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=48150 $D=0
M1228 369 66 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=43520 $D=0
M1229 370 66 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=48150 $D=0
M1230 371 367 211 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=43520 $D=0
M1231 372 368 212 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=48150 $D=0
M1232 168 371 718 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=43520 $D=0
M1233 169 372 719 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=48150 $D=0
M1234 373 718 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=43520 $D=0
M1235 374 719 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=48150 $D=0
M1236 371 65 373 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=43520 $D=0
M1237 372 65 374 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=48150 $D=0
M1238 373 369 221 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=43520 $D=0
M1239 374 370 222 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=48150 $D=0
M1240 225 375 373 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=43520 $D=0
M1241 226 376 374 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=48150 $D=0
M1242 375 67 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=43520 $D=0
M1243 376 67 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=48150 $D=0
M1244 168 68 377 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=43520 $D=0
M1245 169 68 378 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=48150 $D=0
M1246 379 69 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=43520 $D=0
M1247 380 69 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=48150 $D=0
M1248 381 377 211 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=43520 $D=0
M1249 382 378 212 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=48150 $D=0
M1250 168 381 720 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=43520 $D=0
M1251 169 382 721 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=48150 $D=0
M1252 383 720 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=43520 $D=0
M1253 384 721 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=48150 $D=0
M1254 381 68 383 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=43520 $D=0
M1255 382 68 384 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=48150 $D=0
M1256 383 379 221 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=43520 $D=0
M1257 384 380 222 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=48150 $D=0
M1258 225 385 383 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=43520 $D=0
M1259 226 386 384 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=48150 $D=0
M1260 385 70 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=43520 $D=0
M1261 386 70 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=48150 $D=0
M1262 168 71 387 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=43520 $D=0
M1263 169 71 388 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=48150 $D=0
M1264 389 72 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=43520 $D=0
M1265 390 72 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=48150 $D=0
M1266 391 387 211 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=43520 $D=0
M1267 392 388 212 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=48150 $D=0
M1268 168 391 722 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=43520 $D=0
M1269 169 392 723 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=48150 $D=0
M1270 393 722 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=43520 $D=0
M1271 394 723 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=48150 $D=0
M1272 391 71 393 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=43520 $D=0
M1273 392 71 394 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=48150 $D=0
M1274 393 389 221 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=43520 $D=0
M1275 394 390 222 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=48150 $D=0
M1276 225 395 393 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=43520 $D=0
M1277 226 396 394 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=48150 $D=0
M1278 395 73 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=43520 $D=0
M1279 396 73 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=48150 $D=0
M1280 168 74 397 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=43520 $D=0
M1281 169 74 398 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=48150 $D=0
M1282 399 75 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=43520 $D=0
M1283 400 75 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=48150 $D=0
M1284 401 397 211 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=43520 $D=0
M1285 402 398 212 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=48150 $D=0
M1286 168 401 724 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=43520 $D=0
M1287 169 402 725 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=48150 $D=0
M1288 403 724 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=43520 $D=0
M1289 404 725 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=48150 $D=0
M1290 401 74 403 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=43520 $D=0
M1291 402 74 404 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=48150 $D=0
M1292 403 399 221 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=43520 $D=0
M1293 404 400 222 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=48150 $D=0
M1294 225 405 403 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=43520 $D=0
M1295 226 406 404 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=48150 $D=0
M1296 405 76 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=43520 $D=0
M1297 406 76 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=48150 $D=0
M1298 168 77 407 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=43520 $D=0
M1299 169 77 408 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=48150 $D=0
M1300 409 78 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=43520 $D=0
M1301 410 78 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=48150 $D=0
M1302 411 407 211 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=43520 $D=0
M1303 412 408 212 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=48150 $D=0
M1304 168 411 726 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=43520 $D=0
M1305 169 412 727 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=48150 $D=0
M1306 413 726 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=43520 $D=0
M1307 414 727 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=48150 $D=0
M1308 411 77 413 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=43520 $D=0
M1309 412 77 414 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=48150 $D=0
M1310 413 409 221 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=43520 $D=0
M1311 414 410 222 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=48150 $D=0
M1312 225 415 413 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=43520 $D=0
M1313 226 416 414 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=48150 $D=0
M1314 415 79 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=43520 $D=0
M1315 416 79 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=48150 $D=0
M1316 168 80 417 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=43520 $D=0
M1317 169 80 418 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=48150 $D=0
M1318 419 81 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=43520 $D=0
M1319 420 81 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=48150 $D=0
M1320 421 417 211 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=43520 $D=0
M1321 422 418 212 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=48150 $D=0
M1322 168 421 728 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=43520 $D=0
M1323 169 422 729 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=48150 $D=0
M1324 423 728 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=43520 $D=0
M1325 424 729 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=48150 $D=0
M1326 421 80 423 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=43520 $D=0
M1327 422 80 424 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=48150 $D=0
M1328 423 419 221 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=43520 $D=0
M1329 424 420 222 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=48150 $D=0
M1330 225 425 423 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=43520 $D=0
M1331 226 426 424 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=48150 $D=0
M1332 425 82 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=43520 $D=0
M1333 426 82 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=48150 $D=0
M1334 168 83 427 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=43520 $D=0
M1335 169 83 428 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=48150 $D=0
M1336 429 84 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=43520 $D=0
M1337 430 84 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=48150 $D=0
M1338 431 427 211 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=43520 $D=0
M1339 432 428 212 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=48150 $D=0
M1340 168 431 730 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=43520 $D=0
M1341 169 432 731 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=48150 $D=0
M1342 433 730 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=43520 $D=0
M1343 434 731 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=48150 $D=0
M1344 431 83 433 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=43520 $D=0
M1345 432 83 434 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=48150 $D=0
M1346 433 429 221 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=43520 $D=0
M1347 434 430 222 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=48150 $D=0
M1348 225 435 433 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=43520 $D=0
M1349 226 436 434 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=48150 $D=0
M1350 435 85 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=43520 $D=0
M1351 436 85 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=48150 $D=0
M1352 168 86 437 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=43520 $D=0
M1353 169 86 438 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=48150 $D=0
M1354 439 87 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=43520 $D=0
M1355 440 87 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=48150 $D=0
M1356 441 437 211 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=43520 $D=0
M1357 442 438 212 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=48150 $D=0
M1358 168 441 732 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=43520 $D=0
M1359 169 442 733 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=48150 $D=0
M1360 443 732 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=43520 $D=0
M1361 444 733 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=48150 $D=0
M1362 441 86 443 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=43520 $D=0
M1363 442 86 444 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=48150 $D=0
M1364 443 439 221 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=43520 $D=0
M1365 444 440 222 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=48150 $D=0
M1366 225 445 443 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=43520 $D=0
M1367 226 446 444 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=48150 $D=0
M1368 445 88 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=43520 $D=0
M1369 446 88 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=48150 $D=0
M1370 168 89 447 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=43520 $D=0
M1371 169 89 448 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=48150 $D=0
M1372 449 90 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=43520 $D=0
M1373 450 90 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=48150 $D=0
M1374 451 447 211 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=43520 $D=0
M1375 452 448 212 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=48150 $D=0
M1376 168 451 734 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=43520 $D=0
M1377 169 452 735 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=48150 $D=0
M1378 453 734 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=43520 $D=0
M1379 454 735 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=48150 $D=0
M1380 451 89 453 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=43520 $D=0
M1381 452 89 454 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=48150 $D=0
M1382 453 449 221 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=43520 $D=0
M1383 454 450 222 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=48150 $D=0
M1384 225 455 453 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=43520 $D=0
M1385 226 456 454 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=48150 $D=0
M1386 455 91 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=43520 $D=0
M1387 456 91 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=48150 $D=0
M1388 168 92 457 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=43520 $D=0
M1389 169 92 458 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=48150 $D=0
M1390 459 93 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=43520 $D=0
M1391 460 93 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=48150 $D=0
M1392 461 457 211 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=43520 $D=0
M1393 462 458 212 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=48150 $D=0
M1394 168 461 736 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=43520 $D=0
M1395 169 462 737 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=48150 $D=0
M1396 463 736 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=43520 $D=0
M1397 464 737 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=48150 $D=0
M1398 461 92 463 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=43520 $D=0
M1399 462 92 464 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=48150 $D=0
M1400 463 459 221 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=43520 $D=0
M1401 464 460 222 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=48150 $D=0
M1402 225 465 463 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=43520 $D=0
M1403 226 466 464 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=48150 $D=0
M1404 465 94 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=43520 $D=0
M1405 466 94 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=48150 $D=0
M1406 168 95 467 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=43520 $D=0
M1407 169 95 468 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=48150 $D=0
M1408 469 96 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=43520 $D=0
M1409 470 96 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=48150 $D=0
M1410 471 467 211 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=43520 $D=0
M1411 472 468 212 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=48150 $D=0
M1412 168 471 738 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=43520 $D=0
M1413 169 472 739 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=48150 $D=0
M1414 473 738 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=43520 $D=0
M1415 474 739 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=48150 $D=0
M1416 471 95 473 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=43520 $D=0
M1417 472 95 474 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=48150 $D=0
M1418 473 469 221 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=43520 $D=0
M1419 474 470 222 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=48150 $D=0
M1420 225 475 473 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=43520 $D=0
M1421 226 476 474 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=48150 $D=0
M1422 475 97 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=43520 $D=0
M1423 476 97 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=48150 $D=0
M1424 168 98 477 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=43520 $D=0
M1425 169 98 478 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=48150 $D=0
M1426 479 99 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=43520 $D=0
M1427 480 99 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=48150 $D=0
M1428 481 477 211 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=43520 $D=0
M1429 482 478 212 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=48150 $D=0
M1430 168 481 740 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=43520 $D=0
M1431 169 482 741 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=48150 $D=0
M1432 483 740 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=43520 $D=0
M1433 484 741 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=48150 $D=0
M1434 481 98 483 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=43520 $D=0
M1435 482 98 484 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=48150 $D=0
M1436 483 479 221 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=43520 $D=0
M1437 484 480 222 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=48150 $D=0
M1438 225 485 483 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=43520 $D=0
M1439 226 486 484 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=48150 $D=0
M1440 485 100 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=43520 $D=0
M1441 486 100 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=48150 $D=0
M1442 168 101 487 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=43520 $D=0
M1443 169 101 488 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=48150 $D=0
M1444 489 102 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=43520 $D=0
M1445 490 102 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=48150 $D=0
M1446 491 487 211 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=43520 $D=0
M1447 492 488 212 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=48150 $D=0
M1448 168 491 742 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=43520 $D=0
M1449 169 492 743 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=48150 $D=0
M1450 493 742 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=43520 $D=0
M1451 494 743 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=48150 $D=0
M1452 491 101 493 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=43520 $D=0
M1453 492 101 494 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=48150 $D=0
M1454 493 489 221 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=43520 $D=0
M1455 494 490 222 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=48150 $D=0
M1456 225 495 493 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=43520 $D=0
M1457 226 496 494 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=48150 $D=0
M1458 495 103 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=43520 $D=0
M1459 496 103 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=48150 $D=0
M1460 168 104 497 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=43520 $D=0
M1461 169 104 498 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=48150 $D=0
M1462 499 105 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=43520 $D=0
M1463 500 105 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=48150 $D=0
M1464 501 497 211 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=43520 $D=0
M1465 502 498 212 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=48150 $D=0
M1466 168 501 744 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=43520 $D=0
M1467 169 502 745 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=48150 $D=0
M1468 503 744 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=43520 $D=0
M1469 504 745 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=48150 $D=0
M1470 501 104 503 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=43520 $D=0
M1471 502 104 504 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=48150 $D=0
M1472 503 499 221 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=43520 $D=0
M1473 504 500 222 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=48150 $D=0
M1474 225 505 503 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=43520 $D=0
M1475 226 506 504 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=48150 $D=0
M1476 505 106 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=43520 $D=0
M1477 506 106 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=48150 $D=0
M1478 168 107 507 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=43520 $D=0
M1479 169 107 508 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=48150 $D=0
M1480 509 108 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=43520 $D=0
M1481 510 108 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=48150 $D=0
M1482 511 507 211 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=43520 $D=0
M1483 512 508 212 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=48150 $D=0
M1484 168 511 746 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=43520 $D=0
M1485 169 512 747 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=48150 $D=0
M1486 513 746 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=43520 $D=0
M1487 514 747 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=48150 $D=0
M1488 511 107 513 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=43520 $D=0
M1489 512 107 514 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=48150 $D=0
M1490 513 509 221 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=43520 $D=0
M1491 514 510 222 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=48150 $D=0
M1492 225 515 513 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=43520 $D=0
M1493 226 516 514 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=48150 $D=0
M1494 515 109 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=43520 $D=0
M1495 516 109 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=48150 $D=0
M1496 168 110 517 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=43520 $D=0
M1497 169 110 518 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=48150 $D=0
M1498 519 111 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=43520 $D=0
M1499 520 111 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=48150 $D=0
M1500 521 517 211 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=43520 $D=0
M1501 522 518 212 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=48150 $D=0
M1502 168 521 748 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=43520 $D=0
M1503 169 522 749 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=48150 $D=0
M1504 523 748 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=43520 $D=0
M1505 524 749 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=48150 $D=0
M1506 521 110 523 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=43520 $D=0
M1507 522 110 524 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=48150 $D=0
M1508 523 519 221 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=43520 $D=0
M1509 524 520 222 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=48150 $D=0
M1510 225 525 523 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=43520 $D=0
M1511 226 526 524 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=48150 $D=0
M1512 525 112 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=43520 $D=0
M1513 526 112 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=48150 $D=0
M1514 168 113 527 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=43520 $D=0
M1515 169 113 528 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=48150 $D=0
M1516 529 114 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=43520 $D=0
M1517 530 114 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=48150 $D=0
M1518 6 529 221 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=43520 $D=0
M1519 7 530 222 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=48150 $D=0
M1520 225 527 6 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=43520 $D=0
M1521 226 528 7 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=48150 $D=0
M1522 168 533 531 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=43520 $D=0
M1523 169 534 532 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=48150 $D=0
M1524 533 115 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=43520 $D=0
M1525 534 115 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=48150 $D=0
M1526 750 221 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=43520 $D=0
M1527 751 222 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=48150 $D=0
M1528 535 533 750 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=43520 $D=0
M1529 536 534 751 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=48150 $D=0
M1530 168 535 537 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=43520 $D=0
M1531 169 536 538 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=48150 $D=0
M1532 752 537 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=43520 $D=0
M1533 753 538 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=48150 $D=0
M1534 535 531 752 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=43520 $D=0
M1535 536 532 753 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=48150 $D=0
M1536 168 541 539 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=43520 $D=0
M1537 169 542 540 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=48150 $D=0
M1538 541 115 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=43520 $D=0
M1539 542 115 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=48150 $D=0
M1540 754 225 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=43520 $D=0
M1541 755 226 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=48150 $D=0
M1542 543 541 754 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=43520 $D=0
M1543 544 542 755 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=48150 $D=0
M1544 168 543 116 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=43520 $D=0
M1545 169 544 117 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=48150 $D=0
M1546 756 116 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=43520 $D=0
M1547 757 117 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=48150 $D=0
M1548 543 539 756 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=43520 $D=0
M1549 544 540 757 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=48150 $D=0
M1550 545 118 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=43520 $D=0
M1551 546 118 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=48150 $D=0
M1552 547 118 537 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=43520 $D=0
M1553 548 118 538 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=48150 $D=0
M1554 119 545 547 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=43520 $D=0
M1555 120 546 548 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=48150 $D=0
M1556 549 121 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=43520 $D=0
M1557 550 121 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=48150 $D=0
M1558 551 121 116 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=43520 $D=0
M1559 552 121 117 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=48150 $D=0
M1560 758 549 551 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=43520 $D=0
M1561 759 550 552 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=48150 $D=0
M1562 168 116 758 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=43520 $D=0
M1563 169 117 759 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=48150 $D=0
M1564 553 122 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=43520 $D=0
M1565 554 122 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=48150 $D=0
M1566 555 122 551 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=43520 $D=0
M1567 556 122 552 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=48150 $D=0
M1568 12 553 555 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=43520 $D=0
M1569 13 554 556 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=48150 $D=0
M1570 559 557 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=43520 $D=0
M1571 560 558 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=48150 $D=0
M1572 168 563 561 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=43520 $D=0
M1573 169 564 562 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=48150 $D=0
M1574 565 547 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=43520 $D=0
M1575 566 548 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=48150 $D=0
M1576 563 547 557 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=43520 $D=0
M1577 564 548 558 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=48150 $D=0
M1578 559 565 563 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=43520 $D=0
M1579 560 566 564 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=48150 $D=0
M1580 567 561 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=43520 $D=0
M1581 568 562 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=48150 $D=0
M1582 123 561 555 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=43520 $D=0
M1583 557 562 556 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=48150 $D=0
M1584 547 567 123 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=43520 $D=0
M1585 548 568 557 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=48150 $D=0
M1586 569 123 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=43520 $D=0
M1587 570 557 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=48150 $D=0
M1588 571 561 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=43520 $D=0
M1589 572 562 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=48150 $D=0
M1590 573 561 569 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=43520 $D=0
M1591 574 562 570 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=48150 $D=0
M1592 555 571 573 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=43520 $D=0
M1593 556 572 574 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=48150 $D=0
M1594 778 547 168 168 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=43160 $D=0
M1595 779 548 169 169 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=47790 $D=0
M1596 575 555 778 168 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=43160 $D=0
M1597 576 556 779 169 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=47790 $D=0
M1598 577 573 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=43520 $D=0
M1599 578 574 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=48150 $D=0
M1600 579 547 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=43520 $D=0
M1601 580 548 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=48150 $D=0
M1602 168 555 579 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=43520 $D=0
M1603 169 556 580 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=48150 $D=0
M1604 581 547 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=43520 $D=0
M1605 582 548 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=48150 $D=0
M1606 168 555 581 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=43520 $D=0
M1607 169 556 582 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=48150 $D=0
M1608 780 547 168 168 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=43340 $D=0
M1609 781 548 169 169 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=47970 $D=0
M1610 585 555 780 168 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=43340 $D=0
M1611 586 556 781 169 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=47970 $D=0
M1612 168 581 585 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=43520 $D=0
M1613 169 582 586 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=48150 $D=0
M1614 587 128 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=43520 $D=0
M1615 588 128 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=48150 $D=0
M1616 589 128 575 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=43520 $D=0
M1617 590 128 576 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=48150 $D=0
M1618 579 587 589 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=43520 $D=0
M1619 580 588 590 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=48150 $D=0
M1620 591 128 577 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=43520 $D=0
M1621 592 128 578 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=48150 $D=0
M1622 585 587 591 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=43520 $D=0
M1623 586 588 592 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=48150 $D=0
M1624 593 129 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=43520 $D=0
M1625 594 129 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=48150 $D=0
M1626 595 129 591 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=43520 $D=0
M1627 596 129 592 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=48150 $D=0
M1628 589 593 595 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=43520 $D=0
M1629 590 594 596 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=48150 $D=0
M1630 14 595 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=43520 $D=0
M1631 15 596 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=48150 $D=0
M1632 597 130 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=43520 $D=0
M1633 598 130 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=48150 $D=0
M1634 599 130 131 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=43520 $D=0
M1635 600 130 132 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=48150 $D=0
M1636 133 597 599 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=43520 $D=0
M1637 134 598 600 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=48150 $D=0
M1638 601 130 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=43520 $D=0
M1639 602 130 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=48150 $D=0
M1640 604 130 135 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=43520 $D=0
M1641 605 130 137 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=48150 $D=0
M1642 138 601 604 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=43520 $D=0
M1643 136 602 605 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=48150 $D=0
M1644 606 130 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=43520 $D=0
M1645 607 130 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=48150 $D=0
M1646 608 130 127 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=43520 $D=0
M1647 609 130 126 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=48150 $D=0
M1648 139 606 608 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=43520 $D=0
M1649 140 607 609 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=48150 $D=0
M1650 610 130 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=43520 $D=0
M1651 611 130 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=48150 $D=0
M1652 612 130 141 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=43520 $D=0
M1653 613 130 142 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=48150 $D=0
M1654 143 610 612 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=43520 $D=0
M1655 144 611 613 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=48150 $D=0
M1656 614 130 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=43520 $D=0
M1657 615 130 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=48150 $D=0
M1658 616 130 145 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=43520 $D=0
M1659 617 130 146 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=48150 $D=0
M1660 147 614 616 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=43520 $D=0
M1661 147 615 617 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=48150 $D=0
M1662 168 547 768 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=43520 $D=0
M1663 169 548 769 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=48150 $D=0
M1664 134 768 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=43520 $D=0
M1665 131 769 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=48150 $D=0
M1666 618 148 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=43520 $D=0
M1667 619 148 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=48150 $D=0
M1668 149 148 134 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=43520 $D=0
M1669 150 148 131 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=48150 $D=0
M1670 599 618 149 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=43520 $D=0
M1671 600 619 150 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=48150 $D=0
M1672 620 151 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=43520 $D=0
M1673 621 151 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=48150 $D=0
M1674 152 151 149 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=43520 $D=0
M1675 125 151 150 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=48150 $D=0
M1676 604 620 152 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=43520 $D=0
M1677 605 621 125 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=48150 $D=0
M1678 622 153 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=43520 $D=0
M1679 623 153 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=48150 $D=0
M1680 154 153 152 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=43520 $D=0
M1681 155 153 125 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=48150 $D=0
M1682 608 622 154 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=43520 $D=0
M1683 609 623 155 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=48150 $D=0
M1684 624 156 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=43520 $D=0
M1685 625 156 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=48150 $D=0
M1686 157 156 154 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=43520 $D=0
M1687 158 156 155 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=48150 $D=0
M1688 612 624 157 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=43520 $D=0
M1689 613 625 158 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=48150 $D=0
M1690 626 159 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=43520 $D=0
M1691 627 159 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=48150 $D=0
M1692 16 159 157 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=43520 $D=0
M1693 17 159 158 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=48150 $D=0
M1694 616 626 16 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=43520 $D=0
M1695 617 627 17 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=48150 $D=0
M1696 628 160 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=43520 $D=0
M1697 629 160 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=48150 $D=0
M1698 630 160 116 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=43520 $D=0
M1699 631 160 117 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=48150 $D=0
M1700 12 628 630 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=43520 $D=0
M1701 13 629 631 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=48150 $D=0
M1702 632 537 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=43520 $D=0
M1703 633 538 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=48150 $D=0
M1704 168 630 632 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=43520 $D=0
M1705 169 631 633 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=48150 $D=0
M1706 782 537 168 168 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=43340 $D=0
M1707 783 538 169 169 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=47970 $D=0
M1708 636 630 782 168 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=43340 $D=0
M1709 637 631 783 169 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=47970 $D=0
M1710 168 632 636 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=43520 $D=0
M1711 169 633 637 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=48150 $D=0
M1712 770 161 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=43520 $D=0
M1713 771 638 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=48150 $D=0
M1714 168 636 770 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=43520 $D=0
M1715 169 637 771 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=48150 $D=0
M1716 638 770 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=43520 $D=0
M1717 639 771 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=48150 $D=0
M1718 784 537 168 168 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=43160 $D=0
M1719 785 538 169 169 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=47790 $D=0
M1720 640 642 784 168 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=43160 $D=0
M1721 641 643 785 169 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=47790 $D=0
M1722 642 630 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=43520 $D=0
M1723 643 631 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=48150 $D=0
M1724 644 640 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=43520 $D=0
M1725 645 641 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=48150 $D=0
M1726 168 161 644 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=43520 $D=0
M1727 169 638 645 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=48150 $D=0
M1728 647 162 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=43520 $D=0
M1729 648 646 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=48150 $D=0
M1730 646 644 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=43520 $D=0
M1731 163 645 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=48150 $D=0
M1732 168 647 646 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=43520 $D=0
M1733 169 648 163 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=48150 $D=0
M1734 650 649 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=43520 $D=0
M1735 651 164 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=48150 $D=0
M1736 168 654 652 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=43520 $D=0
M1737 169 655 653 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=48150 $D=0
M1738 656 119 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=43520 $D=0
M1739 657 120 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=48150 $D=0
M1740 654 119 649 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=43520 $D=0
M1741 655 120 164 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=48150 $D=0
M1742 650 656 654 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=43520 $D=0
M1743 651 657 655 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=48150 $D=0
M1744 658 652 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=43520 $D=0
M1745 659 653 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=48150 $D=0
M1746 165 652 6 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=43520 $D=0
M1747 649 653 7 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=48150 $D=0
M1748 119 658 165 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=43520 $D=0
M1749 120 659 649 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=48150 $D=0
M1750 660 165 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=43520 $D=0
M1751 661 649 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=48150 $D=0
M1752 662 652 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=43520 $D=0
M1753 663 653 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=48150 $D=0
M1754 199 652 660 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=43520 $D=0
M1755 200 653 661 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=48150 $D=0
M1756 6 662 199 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=43520 $D=0
M1757 7 663 200 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=48150 $D=0
M1758 664 166 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=43520 $D=0
M1759 665 166 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=48150 $D=0
M1760 666 166 199 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=43520 $D=0
M1761 667 166 200 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=48150 $D=0
M1762 14 664 666 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=43520 $D=0
M1763 15 665 667 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=48150 $D=0
M1764 668 167 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=43520 $D=0
M1765 669 167 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=48150 $D=0
M1766 167 167 666 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=43520 $D=0
M1767 167 167 667 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=48150 $D=0
M1768 6 668 167 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=43520 $D=0
M1769 7 669 167 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=48150 $D=0
M1770 670 115 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=43520 $D=0
M1771 671 115 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=48150 $D=0
M1772 168 670 672 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=43520 $D=0
M1773 169 671 673 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=48150 $D=0
M1774 674 115 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=43520 $D=0
M1775 675 115 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=48150 $D=0
M1776 676 672 167 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=43520 $D=0
M1777 677 673 167 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=48150 $D=0
M1778 168 676 772 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=43520 $D=0
M1779 169 677 773 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=48150 $D=0
M1780 678 772 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=43520 $D=0
M1781 679 773 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=48150 $D=0
M1782 676 670 678 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=43520 $D=0
M1783 677 671 679 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=48150 $D=0
M1784 680 674 678 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=43520 $D=0
M1785 681 675 679 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=48150 $D=0
M1786 168 684 682 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=43520 $D=0
M1787 169 685 683 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=48150 $D=0
M1788 684 115 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=43520 $D=0
M1789 685 115 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=48150 $D=0
M1790 774 680 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=43520 $D=0
M1791 775 681 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=48150 $D=0
M1792 686 684 774 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=43520 $D=0
M1793 687 685 775 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=48150 $D=0
M1794 168 686 119 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=43520 $D=0
M1795 169 687 120 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=48150 $D=0
M1796 776 119 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=43520 $D=0
M1797 777 120 169 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=48150 $D=0
M1798 686 682 776 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=43520 $D=0
M1799 687 683 777 169 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=48150 $D=0
.ENDS
***************************************
.SUBCKT ICV_38 1 2 3 4 5 6 7 9 10 11 12 13 14 15 16 17 18 19 20 21
+ 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41
+ 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61
+ 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81
+ 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101
+ 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121
+ 122 123 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141 142
+ 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162
+ 163 164 165 166 167 168
** N=794 EP=166 IP=1514 FDC=1800
M0 172 1 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=33010 $D=1
M1 173 1 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=37640 $D=1
M2 174 172 2 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=33010 $D=1
M3 175 173 3 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=37640 $D=1
M4 6 1 174 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=33010 $D=1
M5 7 1 175 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=37640 $D=1
M6 176 172 4 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=33010 $D=1
M7 177 173 4 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=37640 $D=1
M8 5 1 176 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=33010 $D=1
M9 5 1 177 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=37640 $D=1
M10 178 172 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=33010 $D=1
M11 179 173 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=37640 $D=1
M12 6 1 178 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=33010 $D=1
M13 7 1 179 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=37640 $D=1
M14 182 180 178 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=33010 $D=1
M15 183 181 179 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=37640 $D=1
M16 180 9 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=33010 $D=1
M17 181 9 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=37640 $D=1
M18 184 180 176 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=33010 $D=1
M19 185 181 177 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=37640 $D=1
M20 174 9 184 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=33010 $D=1
M21 175 9 185 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=37640 $D=1
M22 186 10 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=33010 $D=1
M23 187 10 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=37640 $D=1
M24 188 186 184 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=33010 $D=1
M25 189 187 185 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=37640 $D=1
M26 182 10 188 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=33010 $D=1
M27 183 10 189 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=37640 $D=1
M28 190 11 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=33010 $D=1
M29 191 11 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=37640 $D=1
M30 192 190 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=33010 $D=1
M31 193 191 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=37640 $D=1
M32 12 11 192 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=33010 $D=1
M33 13 11 193 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=37640 $D=1
M34 194 190 14 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=33010 $D=1
M35 195 191 15 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=37640 $D=1
M36 196 11 194 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=33010 $D=1
M37 197 11 195 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=37640 $D=1
M38 200 190 198 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=33010 $D=1
M39 201 191 199 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=37640 $D=1
M40 188 11 200 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=33010 $D=1
M41 189 11 201 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=37640 $D=1
M42 204 202 200 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=33010 $D=1
M43 205 203 201 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=37640 $D=1
M44 202 16 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=33010 $D=1
M45 203 16 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=37640 $D=1
M46 206 202 194 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=33010 $D=1
M47 207 203 195 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=37640 $D=1
M48 192 16 206 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=33010 $D=1
M49 193 16 207 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=37640 $D=1
M50 208 17 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=33010 $D=1
M51 209 17 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=37640 $D=1
M52 210 208 206 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=33010 $D=1
M53 211 209 207 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=37640 $D=1
M54 204 17 210 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=33010 $D=1
M55 205 17 211 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=37640 $D=1
M56 6 18 212 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=33010 $D=1
M57 7 18 213 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=37640 $D=1
M58 214 19 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=33010 $D=1
M59 215 19 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=37640 $D=1
M60 216 18 210 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=33010 $D=1
M61 217 18 211 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=37640 $D=1
M62 6 216 685 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=33010 $D=1
M63 7 217 686 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=37640 $D=1
M64 218 685 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=33010 $D=1
M65 219 686 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=37640 $D=1
M66 216 212 218 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=33010 $D=1
M67 217 213 219 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=37640 $D=1
M68 218 19 220 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=33010 $D=1
M69 219 19 221 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=37640 $D=1
M70 224 20 218 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=33010 $D=1
M71 225 20 219 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=37640 $D=1
M72 222 20 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=33010 $D=1
M73 223 20 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=37640 $D=1
M74 6 21 226 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=33010 $D=1
M75 7 21 227 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=37640 $D=1
M76 228 22 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=33010 $D=1
M77 229 22 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=37640 $D=1
M78 230 21 210 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=33010 $D=1
M79 231 21 211 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=37640 $D=1
M80 6 230 687 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=33010 $D=1
M81 7 231 688 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=37640 $D=1
M82 232 687 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=33010 $D=1
M83 233 688 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=37640 $D=1
M84 230 226 232 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=33010 $D=1
M85 231 227 233 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=37640 $D=1
M86 232 22 220 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=33010 $D=1
M87 233 22 221 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=37640 $D=1
M88 224 23 232 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=33010 $D=1
M89 225 23 233 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=37640 $D=1
M90 234 23 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=33010 $D=1
M91 235 23 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=37640 $D=1
M92 6 24 236 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=33010 $D=1
M93 7 24 237 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=37640 $D=1
M94 238 25 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=33010 $D=1
M95 239 25 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=37640 $D=1
M96 240 24 210 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=33010 $D=1
M97 241 24 211 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=37640 $D=1
M98 6 240 689 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=33010 $D=1
M99 7 241 690 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=37640 $D=1
M100 242 689 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=33010 $D=1
M101 243 690 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=37640 $D=1
M102 240 236 242 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=33010 $D=1
M103 241 237 243 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=37640 $D=1
M104 242 25 220 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=33010 $D=1
M105 243 25 221 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=37640 $D=1
M106 224 26 242 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=33010 $D=1
M107 225 26 243 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=37640 $D=1
M108 244 26 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=33010 $D=1
M109 245 26 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=37640 $D=1
M110 6 27 246 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=33010 $D=1
M111 7 27 247 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=37640 $D=1
M112 248 28 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=33010 $D=1
M113 249 28 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=37640 $D=1
M114 250 27 210 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=33010 $D=1
M115 251 27 211 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=37640 $D=1
M116 6 250 691 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=33010 $D=1
M117 7 251 692 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=37640 $D=1
M118 252 691 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=33010 $D=1
M119 253 692 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=37640 $D=1
M120 250 246 252 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=33010 $D=1
M121 251 247 253 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=37640 $D=1
M122 252 28 220 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=33010 $D=1
M123 253 28 221 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=37640 $D=1
M124 224 29 252 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=33010 $D=1
M125 225 29 253 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=37640 $D=1
M126 254 29 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=33010 $D=1
M127 255 29 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=37640 $D=1
M128 6 30 256 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=33010 $D=1
M129 7 30 257 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=37640 $D=1
M130 258 31 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=33010 $D=1
M131 259 31 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=37640 $D=1
M132 260 30 210 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=33010 $D=1
M133 261 30 211 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=37640 $D=1
M134 6 260 693 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=33010 $D=1
M135 7 261 694 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=37640 $D=1
M136 262 693 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=33010 $D=1
M137 263 694 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=37640 $D=1
M138 260 256 262 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=33010 $D=1
M139 261 257 263 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=37640 $D=1
M140 262 31 220 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=33010 $D=1
M141 263 31 221 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=37640 $D=1
M142 224 32 262 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=33010 $D=1
M143 225 32 263 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=37640 $D=1
M144 264 32 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=33010 $D=1
M145 265 32 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=37640 $D=1
M146 6 33 266 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=33010 $D=1
M147 7 33 267 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=37640 $D=1
M148 268 34 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=33010 $D=1
M149 269 34 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=37640 $D=1
M150 270 33 210 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=33010 $D=1
M151 271 33 211 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=37640 $D=1
M152 6 270 695 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=33010 $D=1
M153 7 271 696 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=37640 $D=1
M154 272 695 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=33010 $D=1
M155 273 696 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=37640 $D=1
M156 270 266 272 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=33010 $D=1
M157 271 267 273 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=37640 $D=1
M158 272 34 220 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=33010 $D=1
M159 273 34 221 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=37640 $D=1
M160 224 35 272 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=33010 $D=1
M161 225 35 273 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=37640 $D=1
M162 274 35 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=33010 $D=1
M163 275 35 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=37640 $D=1
M164 6 36 276 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=33010 $D=1
M165 7 36 277 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=37640 $D=1
M166 278 37 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=33010 $D=1
M167 279 37 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=37640 $D=1
M168 280 36 210 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=33010 $D=1
M169 281 36 211 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=37640 $D=1
M170 6 280 697 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=33010 $D=1
M171 7 281 698 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=37640 $D=1
M172 282 697 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=33010 $D=1
M173 283 698 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=37640 $D=1
M174 280 276 282 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=33010 $D=1
M175 281 277 283 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=37640 $D=1
M176 282 37 220 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=33010 $D=1
M177 283 37 221 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=37640 $D=1
M178 224 38 282 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=33010 $D=1
M179 225 38 283 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=37640 $D=1
M180 284 38 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=33010 $D=1
M181 285 38 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=37640 $D=1
M182 6 39 286 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=33010 $D=1
M183 7 39 287 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=37640 $D=1
M184 288 40 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=33010 $D=1
M185 289 40 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=37640 $D=1
M186 290 39 210 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=33010 $D=1
M187 291 39 211 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=37640 $D=1
M188 6 290 699 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=33010 $D=1
M189 7 291 700 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=37640 $D=1
M190 292 699 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=33010 $D=1
M191 293 700 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=37640 $D=1
M192 290 286 292 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=33010 $D=1
M193 291 287 293 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=37640 $D=1
M194 292 40 220 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=33010 $D=1
M195 293 40 221 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=37640 $D=1
M196 224 41 292 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=33010 $D=1
M197 225 41 293 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=37640 $D=1
M198 294 41 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=33010 $D=1
M199 295 41 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=37640 $D=1
M200 6 42 296 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=33010 $D=1
M201 7 42 297 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=37640 $D=1
M202 298 43 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=33010 $D=1
M203 299 43 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=37640 $D=1
M204 300 42 210 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=33010 $D=1
M205 301 42 211 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=37640 $D=1
M206 6 300 701 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=33010 $D=1
M207 7 301 702 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=37640 $D=1
M208 302 701 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=33010 $D=1
M209 303 702 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=37640 $D=1
M210 300 296 302 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=33010 $D=1
M211 301 297 303 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=37640 $D=1
M212 302 43 220 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=33010 $D=1
M213 303 43 221 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=37640 $D=1
M214 224 44 302 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=33010 $D=1
M215 225 44 303 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=37640 $D=1
M216 304 44 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=33010 $D=1
M217 305 44 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=37640 $D=1
M218 6 45 306 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=33010 $D=1
M219 7 45 307 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=37640 $D=1
M220 308 46 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=33010 $D=1
M221 309 46 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=37640 $D=1
M222 310 45 210 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=33010 $D=1
M223 311 45 211 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=37640 $D=1
M224 6 310 703 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=33010 $D=1
M225 7 311 704 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=37640 $D=1
M226 312 703 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=33010 $D=1
M227 313 704 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=37640 $D=1
M228 310 306 312 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=33010 $D=1
M229 311 307 313 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=37640 $D=1
M230 312 46 220 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=33010 $D=1
M231 313 46 221 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=37640 $D=1
M232 224 47 312 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=33010 $D=1
M233 225 47 313 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=37640 $D=1
M234 314 47 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=33010 $D=1
M235 315 47 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=37640 $D=1
M236 6 48 316 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=33010 $D=1
M237 7 48 317 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=37640 $D=1
M238 318 49 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=33010 $D=1
M239 319 49 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=37640 $D=1
M240 320 48 210 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=33010 $D=1
M241 321 48 211 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=37640 $D=1
M242 6 320 705 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=33010 $D=1
M243 7 321 706 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=37640 $D=1
M244 322 705 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=33010 $D=1
M245 323 706 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=37640 $D=1
M246 320 316 322 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=33010 $D=1
M247 321 317 323 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=37640 $D=1
M248 322 49 220 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=33010 $D=1
M249 323 49 221 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=37640 $D=1
M250 224 50 322 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=33010 $D=1
M251 225 50 323 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=37640 $D=1
M252 324 50 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=33010 $D=1
M253 325 50 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=37640 $D=1
M254 6 51 326 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=33010 $D=1
M255 7 51 327 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=37640 $D=1
M256 328 52 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=33010 $D=1
M257 329 52 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=37640 $D=1
M258 330 51 210 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=33010 $D=1
M259 331 51 211 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=37640 $D=1
M260 6 330 707 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=33010 $D=1
M261 7 331 708 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=37640 $D=1
M262 332 707 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=33010 $D=1
M263 333 708 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=37640 $D=1
M264 330 326 332 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=33010 $D=1
M265 331 327 333 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=37640 $D=1
M266 332 52 220 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=33010 $D=1
M267 333 52 221 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=37640 $D=1
M268 224 53 332 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=33010 $D=1
M269 225 53 333 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=37640 $D=1
M270 334 53 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=33010 $D=1
M271 335 53 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=37640 $D=1
M272 6 54 336 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=33010 $D=1
M273 7 54 337 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=37640 $D=1
M274 338 55 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=33010 $D=1
M275 339 55 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=37640 $D=1
M276 340 54 210 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=33010 $D=1
M277 341 54 211 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=37640 $D=1
M278 6 340 709 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=33010 $D=1
M279 7 341 710 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=37640 $D=1
M280 342 709 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=33010 $D=1
M281 343 710 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=37640 $D=1
M282 340 336 342 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=33010 $D=1
M283 341 337 343 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=37640 $D=1
M284 342 55 220 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=33010 $D=1
M285 343 55 221 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=37640 $D=1
M286 224 56 342 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=33010 $D=1
M287 225 56 343 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=37640 $D=1
M288 344 56 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=33010 $D=1
M289 345 56 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=37640 $D=1
M290 6 57 346 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=33010 $D=1
M291 7 57 347 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=37640 $D=1
M292 348 58 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=33010 $D=1
M293 349 58 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=37640 $D=1
M294 350 57 210 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=33010 $D=1
M295 351 57 211 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=37640 $D=1
M296 6 350 711 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=33010 $D=1
M297 7 351 712 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=37640 $D=1
M298 352 711 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=33010 $D=1
M299 353 712 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=37640 $D=1
M300 350 346 352 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=33010 $D=1
M301 351 347 353 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=37640 $D=1
M302 352 58 220 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=33010 $D=1
M303 353 58 221 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=37640 $D=1
M304 224 59 352 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=33010 $D=1
M305 225 59 353 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=37640 $D=1
M306 354 59 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=33010 $D=1
M307 355 59 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=37640 $D=1
M308 6 60 356 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=33010 $D=1
M309 7 60 357 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=37640 $D=1
M310 358 61 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=33010 $D=1
M311 359 61 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=37640 $D=1
M312 360 60 210 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=33010 $D=1
M313 361 60 211 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=37640 $D=1
M314 6 360 713 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=33010 $D=1
M315 7 361 714 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=37640 $D=1
M316 362 713 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=33010 $D=1
M317 363 714 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=37640 $D=1
M318 360 356 362 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=33010 $D=1
M319 361 357 363 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=37640 $D=1
M320 362 61 220 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=33010 $D=1
M321 363 61 221 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=37640 $D=1
M322 224 62 362 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=33010 $D=1
M323 225 62 363 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=37640 $D=1
M324 364 62 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=33010 $D=1
M325 365 62 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=37640 $D=1
M326 6 63 366 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=33010 $D=1
M327 7 63 367 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=37640 $D=1
M328 368 64 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=33010 $D=1
M329 369 64 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=37640 $D=1
M330 370 63 210 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=33010 $D=1
M331 371 63 211 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=37640 $D=1
M332 6 370 715 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=33010 $D=1
M333 7 371 716 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=37640 $D=1
M334 372 715 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=33010 $D=1
M335 373 716 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=37640 $D=1
M336 370 366 372 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=33010 $D=1
M337 371 367 373 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=37640 $D=1
M338 372 64 220 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=33010 $D=1
M339 373 64 221 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=37640 $D=1
M340 224 65 372 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=33010 $D=1
M341 225 65 373 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=37640 $D=1
M342 374 65 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=33010 $D=1
M343 375 65 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=37640 $D=1
M344 6 66 376 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=33010 $D=1
M345 7 66 377 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=37640 $D=1
M346 378 67 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=33010 $D=1
M347 379 67 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=37640 $D=1
M348 380 66 210 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=33010 $D=1
M349 381 66 211 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=37640 $D=1
M350 6 380 717 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=33010 $D=1
M351 7 381 718 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=37640 $D=1
M352 382 717 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=33010 $D=1
M353 383 718 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=37640 $D=1
M354 380 376 382 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=33010 $D=1
M355 381 377 383 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=37640 $D=1
M356 382 67 220 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=33010 $D=1
M357 383 67 221 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=37640 $D=1
M358 224 68 382 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=33010 $D=1
M359 225 68 383 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=37640 $D=1
M360 384 68 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=33010 $D=1
M361 385 68 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=37640 $D=1
M362 6 69 386 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=33010 $D=1
M363 7 69 387 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=37640 $D=1
M364 388 70 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=33010 $D=1
M365 389 70 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=37640 $D=1
M366 390 69 210 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=33010 $D=1
M367 391 69 211 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=37640 $D=1
M368 6 390 719 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=33010 $D=1
M369 7 391 720 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=37640 $D=1
M370 392 719 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=33010 $D=1
M371 393 720 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=37640 $D=1
M372 390 386 392 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=33010 $D=1
M373 391 387 393 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=37640 $D=1
M374 392 70 220 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=33010 $D=1
M375 393 70 221 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=37640 $D=1
M376 224 71 392 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=33010 $D=1
M377 225 71 393 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=37640 $D=1
M378 394 71 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=33010 $D=1
M379 395 71 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=37640 $D=1
M380 6 72 396 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=33010 $D=1
M381 7 72 397 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=37640 $D=1
M382 398 73 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=33010 $D=1
M383 399 73 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=37640 $D=1
M384 400 72 210 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=33010 $D=1
M385 401 72 211 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=37640 $D=1
M386 6 400 721 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=33010 $D=1
M387 7 401 722 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=37640 $D=1
M388 402 721 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=33010 $D=1
M389 403 722 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=37640 $D=1
M390 400 396 402 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=33010 $D=1
M391 401 397 403 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=37640 $D=1
M392 402 73 220 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=33010 $D=1
M393 403 73 221 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=37640 $D=1
M394 224 74 402 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=33010 $D=1
M395 225 74 403 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=37640 $D=1
M396 404 74 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=33010 $D=1
M397 405 74 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=37640 $D=1
M398 6 75 406 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=33010 $D=1
M399 7 75 407 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=37640 $D=1
M400 408 76 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=33010 $D=1
M401 409 76 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=37640 $D=1
M402 410 75 210 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=33010 $D=1
M403 411 75 211 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=37640 $D=1
M404 6 410 723 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=33010 $D=1
M405 7 411 724 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=37640 $D=1
M406 412 723 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=33010 $D=1
M407 413 724 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=37640 $D=1
M408 410 406 412 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=33010 $D=1
M409 411 407 413 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=37640 $D=1
M410 412 76 220 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=33010 $D=1
M411 413 76 221 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=37640 $D=1
M412 224 77 412 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=33010 $D=1
M413 225 77 413 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=37640 $D=1
M414 414 77 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=33010 $D=1
M415 415 77 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=37640 $D=1
M416 6 78 416 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=33010 $D=1
M417 7 78 417 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=37640 $D=1
M418 418 79 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=33010 $D=1
M419 419 79 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=37640 $D=1
M420 420 78 210 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=33010 $D=1
M421 421 78 211 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=37640 $D=1
M422 6 420 725 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=33010 $D=1
M423 7 421 726 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=37640 $D=1
M424 422 725 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=33010 $D=1
M425 423 726 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=37640 $D=1
M426 420 416 422 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=33010 $D=1
M427 421 417 423 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=37640 $D=1
M428 422 79 220 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=33010 $D=1
M429 423 79 221 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=37640 $D=1
M430 224 80 422 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=33010 $D=1
M431 225 80 423 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=37640 $D=1
M432 424 80 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=33010 $D=1
M433 425 80 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=37640 $D=1
M434 6 81 426 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=33010 $D=1
M435 7 81 427 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=37640 $D=1
M436 428 82 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=33010 $D=1
M437 429 82 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=37640 $D=1
M438 430 81 210 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=33010 $D=1
M439 431 81 211 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=37640 $D=1
M440 6 430 727 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=33010 $D=1
M441 7 431 728 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=37640 $D=1
M442 432 727 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=33010 $D=1
M443 433 728 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=37640 $D=1
M444 430 426 432 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=33010 $D=1
M445 431 427 433 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=37640 $D=1
M446 432 82 220 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=33010 $D=1
M447 433 82 221 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=37640 $D=1
M448 224 83 432 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=33010 $D=1
M449 225 83 433 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=37640 $D=1
M450 434 83 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=33010 $D=1
M451 435 83 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=37640 $D=1
M452 6 84 436 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=33010 $D=1
M453 7 84 437 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=37640 $D=1
M454 438 85 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=33010 $D=1
M455 439 85 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=37640 $D=1
M456 440 84 210 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=33010 $D=1
M457 441 84 211 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=37640 $D=1
M458 6 440 729 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=33010 $D=1
M459 7 441 730 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=37640 $D=1
M460 442 729 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=33010 $D=1
M461 443 730 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=37640 $D=1
M462 440 436 442 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=33010 $D=1
M463 441 437 443 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=37640 $D=1
M464 442 85 220 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=33010 $D=1
M465 443 85 221 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=37640 $D=1
M466 224 86 442 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=33010 $D=1
M467 225 86 443 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=37640 $D=1
M468 444 86 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=33010 $D=1
M469 445 86 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=37640 $D=1
M470 6 87 446 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=33010 $D=1
M471 7 87 447 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=37640 $D=1
M472 448 88 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=33010 $D=1
M473 449 88 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=37640 $D=1
M474 450 87 210 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=33010 $D=1
M475 451 87 211 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=37640 $D=1
M476 6 450 731 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=33010 $D=1
M477 7 451 732 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=37640 $D=1
M478 452 731 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=33010 $D=1
M479 453 732 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=37640 $D=1
M480 450 446 452 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=33010 $D=1
M481 451 447 453 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=37640 $D=1
M482 452 88 220 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=33010 $D=1
M483 453 88 221 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=37640 $D=1
M484 224 89 452 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=33010 $D=1
M485 225 89 453 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=37640 $D=1
M486 454 89 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=33010 $D=1
M487 455 89 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=37640 $D=1
M488 6 90 456 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=33010 $D=1
M489 7 90 457 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=37640 $D=1
M490 458 91 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=33010 $D=1
M491 459 91 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=37640 $D=1
M492 460 90 210 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=33010 $D=1
M493 461 90 211 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=37640 $D=1
M494 6 460 733 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=33010 $D=1
M495 7 461 734 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=37640 $D=1
M496 462 733 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=33010 $D=1
M497 463 734 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=37640 $D=1
M498 460 456 462 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=33010 $D=1
M499 461 457 463 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=37640 $D=1
M500 462 91 220 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=33010 $D=1
M501 463 91 221 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=37640 $D=1
M502 224 92 462 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=33010 $D=1
M503 225 92 463 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=37640 $D=1
M504 464 92 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=33010 $D=1
M505 465 92 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=37640 $D=1
M506 6 93 466 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=33010 $D=1
M507 7 93 467 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=37640 $D=1
M508 468 94 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=33010 $D=1
M509 469 94 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=37640 $D=1
M510 470 93 210 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=33010 $D=1
M511 471 93 211 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=37640 $D=1
M512 6 470 735 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=33010 $D=1
M513 7 471 736 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=37640 $D=1
M514 472 735 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=33010 $D=1
M515 473 736 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=37640 $D=1
M516 470 466 472 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=33010 $D=1
M517 471 467 473 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=37640 $D=1
M518 472 94 220 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=33010 $D=1
M519 473 94 221 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=37640 $D=1
M520 224 95 472 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=33010 $D=1
M521 225 95 473 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=37640 $D=1
M522 474 95 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=33010 $D=1
M523 475 95 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=37640 $D=1
M524 6 96 476 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=33010 $D=1
M525 7 96 477 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=37640 $D=1
M526 478 97 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=33010 $D=1
M527 479 97 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=37640 $D=1
M528 480 96 210 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=33010 $D=1
M529 481 96 211 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=37640 $D=1
M530 6 480 737 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=33010 $D=1
M531 7 481 738 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=37640 $D=1
M532 482 737 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=33010 $D=1
M533 483 738 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=37640 $D=1
M534 480 476 482 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=33010 $D=1
M535 481 477 483 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=37640 $D=1
M536 482 97 220 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=33010 $D=1
M537 483 97 221 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=37640 $D=1
M538 224 98 482 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=33010 $D=1
M539 225 98 483 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=37640 $D=1
M540 484 98 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=33010 $D=1
M541 485 98 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=37640 $D=1
M542 6 99 486 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=33010 $D=1
M543 7 99 487 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=37640 $D=1
M544 488 100 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=33010 $D=1
M545 489 100 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=37640 $D=1
M546 490 99 210 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=33010 $D=1
M547 491 99 211 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=37640 $D=1
M548 6 490 739 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=33010 $D=1
M549 7 491 740 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=37640 $D=1
M550 492 739 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=33010 $D=1
M551 493 740 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=37640 $D=1
M552 490 486 492 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=33010 $D=1
M553 491 487 493 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=37640 $D=1
M554 492 100 220 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=33010 $D=1
M555 493 100 221 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=37640 $D=1
M556 224 101 492 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=33010 $D=1
M557 225 101 493 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=37640 $D=1
M558 494 101 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=33010 $D=1
M559 495 101 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=37640 $D=1
M560 6 102 496 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=33010 $D=1
M561 7 102 497 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=37640 $D=1
M562 498 103 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=33010 $D=1
M563 499 103 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=37640 $D=1
M564 500 102 210 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=33010 $D=1
M565 501 102 211 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=37640 $D=1
M566 6 500 741 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=33010 $D=1
M567 7 501 742 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=37640 $D=1
M568 502 741 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=33010 $D=1
M569 503 742 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=37640 $D=1
M570 500 496 502 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=33010 $D=1
M571 501 497 503 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=37640 $D=1
M572 502 103 220 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=33010 $D=1
M573 503 103 221 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=37640 $D=1
M574 224 104 502 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=33010 $D=1
M575 225 104 503 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=37640 $D=1
M576 504 104 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=33010 $D=1
M577 505 104 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=37640 $D=1
M578 6 105 506 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=33010 $D=1
M579 7 105 507 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=37640 $D=1
M580 508 106 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=33010 $D=1
M581 509 106 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=37640 $D=1
M582 510 105 210 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=33010 $D=1
M583 511 105 211 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=37640 $D=1
M584 6 510 743 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=33010 $D=1
M585 7 511 744 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=37640 $D=1
M586 512 743 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=33010 $D=1
M587 513 744 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=37640 $D=1
M588 510 506 512 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=33010 $D=1
M589 511 507 513 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=37640 $D=1
M590 512 106 220 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=33010 $D=1
M591 513 106 221 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=37640 $D=1
M592 224 107 512 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=33010 $D=1
M593 225 107 513 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=37640 $D=1
M594 514 107 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=33010 $D=1
M595 515 107 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=37640 $D=1
M596 6 108 516 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=33010 $D=1
M597 7 108 517 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=37640 $D=1
M598 518 109 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=33010 $D=1
M599 519 109 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=37640 $D=1
M600 520 108 210 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=33010 $D=1
M601 521 108 211 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=37640 $D=1
M602 6 520 745 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=33010 $D=1
M603 7 521 746 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=37640 $D=1
M604 522 745 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=33010 $D=1
M605 523 746 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=37640 $D=1
M606 520 516 522 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=33010 $D=1
M607 521 517 523 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=37640 $D=1
M608 522 109 220 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=33010 $D=1
M609 523 109 221 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=37640 $D=1
M610 224 110 522 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=33010 $D=1
M611 225 110 523 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=37640 $D=1
M612 524 110 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=33010 $D=1
M613 525 110 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=37640 $D=1
M614 6 111 526 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=33010 $D=1
M615 7 111 527 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=37640 $D=1
M616 528 112 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=33010 $D=1
M617 529 112 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=37640 $D=1
M618 6 112 220 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=33010 $D=1
M619 7 112 221 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=37640 $D=1
M620 224 111 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=33010 $D=1
M621 225 111 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=37640 $D=1
M622 6 532 530 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=33010 $D=1
M623 7 533 531 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=37640 $D=1
M624 532 113 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=33010 $D=1
M625 533 113 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=37640 $D=1
M626 747 220 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=33010 $D=1
M627 748 221 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=37640 $D=1
M628 534 530 747 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=33010 $D=1
M629 535 531 748 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=37640 $D=1
M630 6 534 536 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=33010 $D=1
M631 7 535 537 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=37640 $D=1
M632 749 536 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=33010 $D=1
M633 750 537 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=37640 $D=1
M634 534 532 749 6 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=33010 $D=1
M635 535 533 750 7 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=37640 $D=1
M636 6 540 538 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=33010 $D=1
M637 7 541 539 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=37640 $D=1
M638 540 113 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=33010 $D=1
M639 541 113 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=37640 $D=1
M640 751 224 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=33010 $D=1
M641 752 225 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=37640 $D=1
M642 542 538 751 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=33010 $D=1
M643 543 539 752 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=37640 $D=1
M644 6 542 114 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=33010 $D=1
M645 7 543 115 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=37640 $D=1
M646 753 114 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=33010 $D=1
M647 754 115 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=37640 $D=1
M648 542 540 753 6 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=33010 $D=1
M649 543 541 754 7 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=37640 $D=1
M650 544 116 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=33010 $D=1
M651 545 116 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=37640 $D=1
M652 546 544 536 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=33010 $D=1
M653 547 545 537 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=37640 $D=1
M654 117 116 546 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=33010 $D=1
M655 118 116 547 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=37640 $D=1
M656 548 119 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=33010 $D=1
M657 549 119 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=37640 $D=1
M658 550 548 114 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=33010 $D=1
M659 551 549 115 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=37640 $D=1
M660 755 119 550 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=33010 $D=1
M661 756 119 551 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=37640 $D=1
M662 6 114 755 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=33010 $D=1
M663 7 115 756 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=37640 $D=1
M664 552 120 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=33010 $D=1
M665 553 120 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=37640 $D=1
M666 554 552 550 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=33010 $D=1
M667 555 553 551 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=37640 $D=1
M668 12 120 554 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=33010 $D=1
M669 13 120 555 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=37640 $D=1
M670 557 556 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=33010 $D=1
M671 558 121 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=37640 $D=1
M672 6 561 559 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=33010 $D=1
M673 7 562 560 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=37640 $D=1
M674 563 546 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=33010 $D=1
M675 564 547 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=37640 $D=1
M676 561 563 556 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=33010 $D=1
M677 562 564 121 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=37640 $D=1
M678 557 546 561 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=33010 $D=1
M679 558 547 562 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=37640 $D=1
M680 565 559 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=33010 $D=1
M681 566 560 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=37640 $D=1
M682 122 565 554 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=33010 $D=1
M683 556 566 555 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=37640 $D=1
M684 546 559 122 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=33010 $D=1
M685 547 560 556 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=37640 $D=1
M686 567 122 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=33010 $D=1
M687 568 556 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=37640 $D=1
M688 569 559 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=33010 $D=1
M689 570 560 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=37640 $D=1
M690 571 569 567 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=33010 $D=1
M691 572 570 568 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=37640 $D=1
M692 554 559 571 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=33010 $D=1
M693 555 560 572 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=37640 $D=1
M694 573 546 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=33010 $D=1
M695 574 547 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=37640 $D=1
M696 6 554 573 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=33010 $D=1
M697 7 555 574 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=37640 $D=1
M698 575 571 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=33010 $D=1
M699 576 572 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=37640 $D=1
M700 783 546 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=33010 $D=1
M701 784 547 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=37640 $D=1
M702 577 554 783 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=33010 $D=1
M703 578 555 784 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=37640 $D=1
M704 785 546 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=33010 $D=1
M705 786 547 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=37640 $D=1
M706 579 554 785 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=33010 $D=1
M707 580 555 786 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=37640 $D=1
M708 583 546 581 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=33010 $D=1
M709 584 547 582 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=37640 $D=1
M710 581 554 583 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=33010 $D=1
M711 582 555 584 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=37640 $D=1
M712 6 579 581 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=33010 $D=1
M713 7 580 582 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=37640 $D=1
M714 585 127 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=33010 $D=1
M715 586 127 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=37640 $D=1
M716 587 585 573 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=33010 $D=1
M717 588 586 574 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=37640 $D=1
M718 577 127 587 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=33010 $D=1
M719 578 127 588 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=37640 $D=1
M720 589 585 575 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=33010 $D=1
M721 590 586 576 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=37640 $D=1
M722 583 127 589 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=33010 $D=1
M723 584 127 590 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=37640 $D=1
M724 591 128 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=33010 $D=1
M725 592 128 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=37640 $D=1
M726 593 591 589 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=33010 $D=1
M727 594 592 590 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=37640 $D=1
M728 587 128 593 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=33010 $D=1
M729 588 128 594 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=37640 $D=1
M730 14 593 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=33010 $D=1
M731 15 594 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=37640 $D=1
M732 595 129 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=33010 $D=1
M733 596 129 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=37640 $D=1
M734 597 595 130 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=33010 $D=1
M735 598 596 131 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=37640 $D=1
M736 132 129 597 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=33010 $D=1
M737 133 129 598 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=37640 $D=1
M738 599 129 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=33010 $D=1
M739 600 129 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=37640 $D=1
M740 602 599 134 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=33010 $D=1
M741 603 600 136 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=37640 $D=1
M742 137 129 602 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=33010 $D=1
M743 135 129 603 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=37640 $D=1
M744 604 129 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=33010 $D=1
M745 605 129 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=37640 $D=1
M746 606 604 123 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=33010 $D=1
M747 607 605 126 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=37640 $D=1
M748 138 129 606 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=33010 $D=1
M749 139 129 607 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=37640 $D=1
M750 608 129 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=33010 $D=1
M751 609 129 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=37640 $D=1
M752 610 608 140 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=33010 $D=1
M753 611 609 141 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=37640 $D=1
M754 142 129 610 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=33010 $D=1
M755 143 129 611 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=37640 $D=1
M756 612 129 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=33010 $D=1
M757 613 129 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=37640 $D=1
M758 614 612 144 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=33010 $D=1
M759 615 613 145 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=37640 $D=1
M760 142 129 614 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=33010 $D=1
M761 142 129 615 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=37640 $D=1
M762 6 546 765 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=33010 $D=1
M763 7 547 766 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=37640 $D=1
M764 133 765 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=33010 $D=1
M765 130 766 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=37640 $D=1
M766 616 146 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=33010 $D=1
M767 617 146 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=37640 $D=1
M768 147 616 133 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=33010 $D=1
M769 148 617 130 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=37640 $D=1
M770 597 146 147 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=33010 $D=1
M771 598 146 148 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=37640 $D=1
M772 618 149 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=33010 $D=1
M773 619 149 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=37640 $D=1
M774 150 618 147 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=33010 $D=1
M775 125 619 148 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=37640 $D=1
M776 602 149 150 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=33010 $D=1
M777 603 149 125 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=37640 $D=1
M778 620 151 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=33010 $D=1
M779 621 151 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=37640 $D=1
M780 152 620 150 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=33010 $D=1
M781 153 621 125 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=37640 $D=1
M782 606 151 152 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=33010 $D=1
M783 607 151 153 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=37640 $D=1
M784 622 154 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=33010 $D=1
M785 623 154 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=37640 $D=1
M786 155 622 152 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=33010 $D=1
M787 156 623 153 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=37640 $D=1
M788 610 154 155 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=33010 $D=1
M789 611 154 156 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=37640 $D=1
M790 624 157 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=33010 $D=1
M791 625 157 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=37640 $D=1
M792 196 624 155 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=33010 $D=1
M793 197 625 156 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=37640 $D=1
M794 614 157 196 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=33010 $D=1
M795 615 157 197 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=37640 $D=1
M796 626 158 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=33010 $D=1
M797 627 158 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=37640 $D=1
M798 628 626 114 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=33010 $D=1
M799 629 627 115 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=37640 $D=1
M800 12 158 628 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=33010 $D=1
M801 13 158 629 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=37640 $D=1
M802 787 536 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=33010 $D=1
M803 788 537 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=37640 $D=1
M804 630 628 787 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=33010 $D=1
M805 631 629 788 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=37640 $D=1
M806 634 536 632 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=33010 $D=1
M807 635 537 633 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=37640 $D=1
M808 632 628 634 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=33010 $D=1
M809 633 629 635 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=37640 $D=1
M810 6 630 632 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=33010 $D=1
M811 7 631 633 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=37640 $D=1
M812 789 159 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=33010 $D=1
M813 790 636 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=37640 $D=1
M814 767 634 789 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=33010 $D=1
M815 768 635 790 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=37640 $D=1
M816 636 767 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=33010 $D=1
M817 160 768 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=37640 $D=1
M818 637 536 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=33010 $D=1
M819 638 537 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=37640 $D=1
M820 6 639 637 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=33010 $D=1
M821 7 640 638 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=37640 $D=1
M822 639 628 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=33010 $D=1
M823 640 629 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=37640 $D=1
M824 791 637 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=33010 $D=1
M825 792 638 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=37640 $D=1
M826 641 159 791 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=33010 $D=1
M827 642 636 792 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=37640 $D=1
M828 644 161 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=33010 $D=1
M829 645 643 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=37640 $D=1
M830 793 641 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=33010 $D=1
M831 794 642 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=37640 $D=1
M832 643 644 793 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=33010 $D=1
M833 162 645 794 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=37640 $D=1
M834 647 646 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=33010 $D=1
M835 648 163 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=37640 $D=1
M836 6 651 649 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=33010 $D=1
M837 7 652 650 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=37640 $D=1
M838 653 117 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=33010 $D=1
M839 654 118 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=37640 $D=1
M840 651 653 646 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=33010 $D=1
M841 652 654 163 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=37640 $D=1
M842 647 117 651 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=33010 $D=1
M843 648 118 652 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=37640 $D=1
M844 655 649 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=33010 $D=1
M845 656 650 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=37640 $D=1
M846 164 655 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=33010 $D=1
M847 646 656 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=37640 $D=1
M848 117 649 164 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=33010 $D=1
M849 118 650 646 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=37640 $D=1
M850 657 164 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=33010 $D=1
M851 658 646 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=37640 $D=1
M852 659 649 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=33010 $D=1
M853 660 650 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=37640 $D=1
M854 198 659 657 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=33010 $D=1
M855 199 660 658 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=37640 $D=1
M856 6 649 198 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=33010 $D=1
M857 7 650 199 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=37640 $D=1
M858 661 165 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=33010 $D=1
M859 662 165 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=37640 $D=1
M860 663 661 198 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=33010 $D=1
M861 664 662 199 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=37640 $D=1
M862 14 165 663 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=33010 $D=1
M863 15 165 664 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=37640 $D=1
M864 665 166 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=33010 $D=1
M865 666 166 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=37640 $D=1
M866 166 665 663 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=33010 $D=1
M867 166 666 664 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=37640 $D=1
M868 6 166 166 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=33010 $D=1
M869 7 166 166 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=37640 $D=1
M870 667 113 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=33010 $D=1
M871 668 113 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=37640 $D=1
M872 6 667 669 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=33010 $D=1
M873 7 668 670 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=37640 $D=1
M874 671 113 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=33010 $D=1
M875 672 113 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=37640 $D=1
M876 673 667 166 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=33010 $D=1
M877 674 668 166 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=37640 $D=1
M878 6 673 769 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=33010 $D=1
M879 7 674 770 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=37640 $D=1
M880 675 769 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=33010 $D=1
M881 676 770 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=37640 $D=1
M882 673 669 675 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=33010 $D=1
M883 674 670 676 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=37640 $D=1
M884 677 113 675 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=33010 $D=1
M885 678 113 676 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=37640 $D=1
M886 6 681 679 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=33010 $D=1
M887 7 682 680 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=37640 $D=1
M888 681 113 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=33010 $D=1
M889 682 113 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=37640 $D=1
M890 771 677 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=33010 $D=1
M891 772 678 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=37640 $D=1
M892 683 679 771 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=33010 $D=1
M893 684 680 772 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=37640 $D=1
M894 6 683 117 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=33010 $D=1
M895 7 684 118 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=37640 $D=1
M896 773 117 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=33010 $D=1
M897 774 118 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=37640 $D=1
M898 683 681 773 6 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=33010 $D=1
M899 684 682 774 7 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=37640 $D=1
M900 172 1 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=34260 $D=0
M901 173 1 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=38890 $D=0
M902 174 1 2 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=34260 $D=0
M903 175 1 3 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=38890 $D=0
M904 6 172 174 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=34260 $D=0
M905 7 173 175 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=38890 $D=0
M906 176 1 4 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=34260 $D=0
M907 177 1 4 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=38890 $D=0
M908 5 172 176 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=34260 $D=0
M909 5 173 177 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=38890 $D=0
M910 178 1 6 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=34260 $D=0
M911 179 1 7 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=38890 $D=0
M912 6 172 178 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=34260 $D=0
M913 7 173 179 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=38890 $D=0
M914 182 9 178 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=34260 $D=0
M915 183 9 179 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=38890 $D=0
M916 180 9 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=34260 $D=0
M917 181 9 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=38890 $D=0
M918 184 9 176 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=34260 $D=0
M919 185 9 177 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=38890 $D=0
M920 174 180 184 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=34260 $D=0
M921 175 181 185 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=38890 $D=0
M922 186 10 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=34260 $D=0
M923 187 10 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=38890 $D=0
M924 188 10 184 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=34260 $D=0
M925 189 10 185 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=38890 $D=0
M926 182 186 188 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=34260 $D=0
M927 183 187 189 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=38890 $D=0
M928 190 11 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=34260 $D=0
M929 191 11 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=38890 $D=0
M930 192 11 6 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=34260 $D=0
M931 193 11 7 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=38890 $D=0
M932 12 190 192 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=34260 $D=0
M933 13 191 193 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=38890 $D=0
M934 194 11 14 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=34260 $D=0
M935 195 11 15 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=38890 $D=0
M936 196 190 194 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=34260 $D=0
M937 197 191 195 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=38890 $D=0
M938 200 11 198 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=34260 $D=0
M939 201 11 199 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=38890 $D=0
M940 188 190 200 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=34260 $D=0
M941 189 191 201 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=38890 $D=0
M942 204 16 200 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=34260 $D=0
M943 205 16 201 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=38890 $D=0
M944 202 16 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=34260 $D=0
M945 203 16 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=38890 $D=0
M946 206 16 194 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=34260 $D=0
M947 207 16 195 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=38890 $D=0
M948 192 202 206 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=34260 $D=0
M949 193 203 207 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=38890 $D=0
M950 208 17 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=34260 $D=0
M951 209 17 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=38890 $D=0
M952 210 17 206 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=34260 $D=0
M953 211 17 207 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=38890 $D=0
M954 204 208 210 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=34260 $D=0
M955 205 209 211 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=38890 $D=0
M956 167 18 212 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=34260 $D=0
M957 168 18 213 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=38890 $D=0
M958 214 19 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=34260 $D=0
M959 215 19 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=38890 $D=0
M960 216 212 210 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=34260 $D=0
M961 217 213 211 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=38890 $D=0
M962 167 216 685 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=34260 $D=0
M963 168 217 686 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=38890 $D=0
M964 218 685 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=34260 $D=0
M965 219 686 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=38890 $D=0
M966 216 18 218 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=34260 $D=0
M967 217 18 219 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=38890 $D=0
M968 218 214 220 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=34260 $D=0
M969 219 215 221 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=38890 $D=0
M970 224 222 218 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=34260 $D=0
M971 225 223 219 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=38890 $D=0
M972 222 20 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=34260 $D=0
M973 223 20 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=38890 $D=0
M974 167 21 226 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=34260 $D=0
M975 168 21 227 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=38890 $D=0
M976 228 22 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=34260 $D=0
M977 229 22 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=38890 $D=0
M978 230 226 210 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=34260 $D=0
M979 231 227 211 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=38890 $D=0
M980 167 230 687 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=34260 $D=0
M981 168 231 688 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=38890 $D=0
M982 232 687 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=34260 $D=0
M983 233 688 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=38890 $D=0
M984 230 21 232 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=34260 $D=0
M985 231 21 233 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=38890 $D=0
M986 232 228 220 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=34260 $D=0
M987 233 229 221 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=38890 $D=0
M988 224 234 232 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=34260 $D=0
M989 225 235 233 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=38890 $D=0
M990 234 23 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=34260 $D=0
M991 235 23 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=38890 $D=0
M992 167 24 236 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=34260 $D=0
M993 168 24 237 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=38890 $D=0
M994 238 25 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=34260 $D=0
M995 239 25 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=38890 $D=0
M996 240 236 210 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=34260 $D=0
M997 241 237 211 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=38890 $D=0
M998 167 240 689 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=34260 $D=0
M999 168 241 690 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=38890 $D=0
M1000 242 689 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=34260 $D=0
M1001 243 690 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=38890 $D=0
M1002 240 24 242 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=34260 $D=0
M1003 241 24 243 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=38890 $D=0
M1004 242 238 220 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=34260 $D=0
M1005 243 239 221 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=38890 $D=0
M1006 224 244 242 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=34260 $D=0
M1007 225 245 243 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=38890 $D=0
M1008 244 26 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=34260 $D=0
M1009 245 26 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=38890 $D=0
M1010 167 27 246 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=34260 $D=0
M1011 168 27 247 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=38890 $D=0
M1012 248 28 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=34260 $D=0
M1013 249 28 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=38890 $D=0
M1014 250 246 210 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=34260 $D=0
M1015 251 247 211 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=38890 $D=0
M1016 167 250 691 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=34260 $D=0
M1017 168 251 692 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=38890 $D=0
M1018 252 691 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=34260 $D=0
M1019 253 692 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=38890 $D=0
M1020 250 27 252 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=34260 $D=0
M1021 251 27 253 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=38890 $D=0
M1022 252 248 220 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=34260 $D=0
M1023 253 249 221 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=38890 $D=0
M1024 224 254 252 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=34260 $D=0
M1025 225 255 253 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=38890 $D=0
M1026 254 29 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=34260 $D=0
M1027 255 29 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=38890 $D=0
M1028 167 30 256 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=34260 $D=0
M1029 168 30 257 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=38890 $D=0
M1030 258 31 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=34260 $D=0
M1031 259 31 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=38890 $D=0
M1032 260 256 210 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=34260 $D=0
M1033 261 257 211 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=38890 $D=0
M1034 167 260 693 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=34260 $D=0
M1035 168 261 694 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=38890 $D=0
M1036 262 693 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=34260 $D=0
M1037 263 694 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=38890 $D=0
M1038 260 30 262 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=34260 $D=0
M1039 261 30 263 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=38890 $D=0
M1040 262 258 220 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=34260 $D=0
M1041 263 259 221 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=38890 $D=0
M1042 224 264 262 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=34260 $D=0
M1043 225 265 263 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=38890 $D=0
M1044 264 32 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=34260 $D=0
M1045 265 32 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=38890 $D=0
M1046 167 33 266 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=34260 $D=0
M1047 168 33 267 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=38890 $D=0
M1048 268 34 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=34260 $D=0
M1049 269 34 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=38890 $D=0
M1050 270 266 210 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=34260 $D=0
M1051 271 267 211 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=38890 $D=0
M1052 167 270 695 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=34260 $D=0
M1053 168 271 696 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=38890 $D=0
M1054 272 695 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=34260 $D=0
M1055 273 696 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=38890 $D=0
M1056 270 33 272 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=34260 $D=0
M1057 271 33 273 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=38890 $D=0
M1058 272 268 220 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=34260 $D=0
M1059 273 269 221 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=38890 $D=0
M1060 224 274 272 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=34260 $D=0
M1061 225 275 273 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=38890 $D=0
M1062 274 35 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=34260 $D=0
M1063 275 35 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=38890 $D=0
M1064 167 36 276 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=34260 $D=0
M1065 168 36 277 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=38890 $D=0
M1066 278 37 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=34260 $D=0
M1067 279 37 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=38890 $D=0
M1068 280 276 210 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=34260 $D=0
M1069 281 277 211 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=38890 $D=0
M1070 167 280 697 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=34260 $D=0
M1071 168 281 698 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=38890 $D=0
M1072 282 697 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=34260 $D=0
M1073 283 698 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=38890 $D=0
M1074 280 36 282 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=34260 $D=0
M1075 281 36 283 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=38890 $D=0
M1076 282 278 220 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=34260 $D=0
M1077 283 279 221 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=38890 $D=0
M1078 224 284 282 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=34260 $D=0
M1079 225 285 283 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=38890 $D=0
M1080 284 38 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=34260 $D=0
M1081 285 38 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=38890 $D=0
M1082 167 39 286 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=34260 $D=0
M1083 168 39 287 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=38890 $D=0
M1084 288 40 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=34260 $D=0
M1085 289 40 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=38890 $D=0
M1086 290 286 210 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=34260 $D=0
M1087 291 287 211 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=38890 $D=0
M1088 167 290 699 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=34260 $D=0
M1089 168 291 700 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=38890 $D=0
M1090 292 699 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=34260 $D=0
M1091 293 700 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=38890 $D=0
M1092 290 39 292 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=34260 $D=0
M1093 291 39 293 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=38890 $D=0
M1094 292 288 220 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=34260 $D=0
M1095 293 289 221 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=38890 $D=0
M1096 224 294 292 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=34260 $D=0
M1097 225 295 293 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=38890 $D=0
M1098 294 41 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=34260 $D=0
M1099 295 41 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=38890 $D=0
M1100 167 42 296 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=34260 $D=0
M1101 168 42 297 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=38890 $D=0
M1102 298 43 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=34260 $D=0
M1103 299 43 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=38890 $D=0
M1104 300 296 210 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=34260 $D=0
M1105 301 297 211 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=38890 $D=0
M1106 167 300 701 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=34260 $D=0
M1107 168 301 702 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=38890 $D=0
M1108 302 701 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=34260 $D=0
M1109 303 702 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=38890 $D=0
M1110 300 42 302 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=34260 $D=0
M1111 301 42 303 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=38890 $D=0
M1112 302 298 220 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=34260 $D=0
M1113 303 299 221 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=38890 $D=0
M1114 224 304 302 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=34260 $D=0
M1115 225 305 303 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=38890 $D=0
M1116 304 44 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=34260 $D=0
M1117 305 44 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=38890 $D=0
M1118 167 45 306 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=34260 $D=0
M1119 168 45 307 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=38890 $D=0
M1120 308 46 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=34260 $D=0
M1121 309 46 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=38890 $D=0
M1122 310 306 210 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=34260 $D=0
M1123 311 307 211 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=38890 $D=0
M1124 167 310 703 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=34260 $D=0
M1125 168 311 704 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=38890 $D=0
M1126 312 703 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=34260 $D=0
M1127 313 704 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=38890 $D=0
M1128 310 45 312 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=34260 $D=0
M1129 311 45 313 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=38890 $D=0
M1130 312 308 220 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=34260 $D=0
M1131 313 309 221 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=38890 $D=0
M1132 224 314 312 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=34260 $D=0
M1133 225 315 313 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=38890 $D=0
M1134 314 47 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=34260 $D=0
M1135 315 47 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=38890 $D=0
M1136 167 48 316 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=34260 $D=0
M1137 168 48 317 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=38890 $D=0
M1138 318 49 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=34260 $D=0
M1139 319 49 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=38890 $D=0
M1140 320 316 210 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=34260 $D=0
M1141 321 317 211 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=38890 $D=0
M1142 167 320 705 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=34260 $D=0
M1143 168 321 706 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=38890 $D=0
M1144 322 705 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=34260 $D=0
M1145 323 706 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=38890 $D=0
M1146 320 48 322 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=34260 $D=0
M1147 321 48 323 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=38890 $D=0
M1148 322 318 220 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=34260 $D=0
M1149 323 319 221 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=38890 $D=0
M1150 224 324 322 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=34260 $D=0
M1151 225 325 323 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=38890 $D=0
M1152 324 50 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=34260 $D=0
M1153 325 50 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=38890 $D=0
M1154 167 51 326 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=34260 $D=0
M1155 168 51 327 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=38890 $D=0
M1156 328 52 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=34260 $D=0
M1157 329 52 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=38890 $D=0
M1158 330 326 210 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=34260 $D=0
M1159 331 327 211 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=38890 $D=0
M1160 167 330 707 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=34260 $D=0
M1161 168 331 708 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=38890 $D=0
M1162 332 707 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=34260 $D=0
M1163 333 708 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=38890 $D=0
M1164 330 51 332 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=34260 $D=0
M1165 331 51 333 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=38890 $D=0
M1166 332 328 220 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=34260 $D=0
M1167 333 329 221 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=38890 $D=0
M1168 224 334 332 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=34260 $D=0
M1169 225 335 333 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=38890 $D=0
M1170 334 53 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=34260 $D=0
M1171 335 53 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=38890 $D=0
M1172 167 54 336 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=34260 $D=0
M1173 168 54 337 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=38890 $D=0
M1174 338 55 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=34260 $D=0
M1175 339 55 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=38890 $D=0
M1176 340 336 210 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=34260 $D=0
M1177 341 337 211 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=38890 $D=0
M1178 167 340 709 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=34260 $D=0
M1179 168 341 710 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=38890 $D=0
M1180 342 709 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=34260 $D=0
M1181 343 710 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=38890 $D=0
M1182 340 54 342 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=34260 $D=0
M1183 341 54 343 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=38890 $D=0
M1184 342 338 220 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=34260 $D=0
M1185 343 339 221 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=38890 $D=0
M1186 224 344 342 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=34260 $D=0
M1187 225 345 343 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=38890 $D=0
M1188 344 56 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=34260 $D=0
M1189 345 56 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=38890 $D=0
M1190 167 57 346 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=34260 $D=0
M1191 168 57 347 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=38890 $D=0
M1192 348 58 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=34260 $D=0
M1193 349 58 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=38890 $D=0
M1194 350 346 210 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=34260 $D=0
M1195 351 347 211 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=38890 $D=0
M1196 167 350 711 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=34260 $D=0
M1197 168 351 712 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=38890 $D=0
M1198 352 711 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=34260 $D=0
M1199 353 712 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=38890 $D=0
M1200 350 57 352 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=34260 $D=0
M1201 351 57 353 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=38890 $D=0
M1202 352 348 220 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=34260 $D=0
M1203 353 349 221 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=38890 $D=0
M1204 224 354 352 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=34260 $D=0
M1205 225 355 353 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=38890 $D=0
M1206 354 59 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=34260 $D=0
M1207 355 59 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=38890 $D=0
M1208 167 60 356 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=34260 $D=0
M1209 168 60 357 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=38890 $D=0
M1210 358 61 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=34260 $D=0
M1211 359 61 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=38890 $D=0
M1212 360 356 210 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=34260 $D=0
M1213 361 357 211 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=38890 $D=0
M1214 167 360 713 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=34260 $D=0
M1215 168 361 714 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=38890 $D=0
M1216 362 713 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=34260 $D=0
M1217 363 714 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=38890 $D=0
M1218 360 60 362 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=34260 $D=0
M1219 361 60 363 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=38890 $D=0
M1220 362 358 220 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=34260 $D=0
M1221 363 359 221 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=38890 $D=0
M1222 224 364 362 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=34260 $D=0
M1223 225 365 363 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=38890 $D=0
M1224 364 62 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=34260 $D=0
M1225 365 62 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=38890 $D=0
M1226 167 63 366 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=34260 $D=0
M1227 168 63 367 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=38890 $D=0
M1228 368 64 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=34260 $D=0
M1229 369 64 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=38890 $D=0
M1230 370 366 210 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=34260 $D=0
M1231 371 367 211 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=38890 $D=0
M1232 167 370 715 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=34260 $D=0
M1233 168 371 716 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=38890 $D=0
M1234 372 715 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=34260 $D=0
M1235 373 716 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=38890 $D=0
M1236 370 63 372 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=34260 $D=0
M1237 371 63 373 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=38890 $D=0
M1238 372 368 220 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=34260 $D=0
M1239 373 369 221 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=38890 $D=0
M1240 224 374 372 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=34260 $D=0
M1241 225 375 373 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=38890 $D=0
M1242 374 65 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=34260 $D=0
M1243 375 65 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=38890 $D=0
M1244 167 66 376 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=34260 $D=0
M1245 168 66 377 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=38890 $D=0
M1246 378 67 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=34260 $D=0
M1247 379 67 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=38890 $D=0
M1248 380 376 210 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=34260 $D=0
M1249 381 377 211 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=38890 $D=0
M1250 167 380 717 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=34260 $D=0
M1251 168 381 718 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=38890 $D=0
M1252 382 717 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=34260 $D=0
M1253 383 718 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=38890 $D=0
M1254 380 66 382 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=34260 $D=0
M1255 381 66 383 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=38890 $D=0
M1256 382 378 220 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=34260 $D=0
M1257 383 379 221 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=38890 $D=0
M1258 224 384 382 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=34260 $D=0
M1259 225 385 383 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=38890 $D=0
M1260 384 68 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=34260 $D=0
M1261 385 68 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=38890 $D=0
M1262 167 69 386 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=34260 $D=0
M1263 168 69 387 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=38890 $D=0
M1264 388 70 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=34260 $D=0
M1265 389 70 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=38890 $D=0
M1266 390 386 210 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=34260 $D=0
M1267 391 387 211 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=38890 $D=0
M1268 167 390 719 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=34260 $D=0
M1269 168 391 720 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=38890 $D=0
M1270 392 719 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=34260 $D=0
M1271 393 720 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=38890 $D=0
M1272 390 69 392 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=34260 $D=0
M1273 391 69 393 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=38890 $D=0
M1274 392 388 220 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=34260 $D=0
M1275 393 389 221 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=38890 $D=0
M1276 224 394 392 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=34260 $D=0
M1277 225 395 393 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=38890 $D=0
M1278 394 71 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=34260 $D=0
M1279 395 71 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=38890 $D=0
M1280 167 72 396 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=34260 $D=0
M1281 168 72 397 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=38890 $D=0
M1282 398 73 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=34260 $D=0
M1283 399 73 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=38890 $D=0
M1284 400 396 210 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=34260 $D=0
M1285 401 397 211 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=38890 $D=0
M1286 167 400 721 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=34260 $D=0
M1287 168 401 722 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=38890 $D=0
M1288 402 721 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=34260 $D=0
M1289 403 722 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=38890 $D=0
M1290 400 72 402 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=34260 $D=0
M1291 401 72 403 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=38890 $D=0
M1292 402 398 220 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=34260 $D=0
M1293 403 399 221 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=38890 $D=0
M1294 224 404 402 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=34260 $D=0
M1295 225 405 403 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=38890 $D=0
M1296 404 74 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=34260 $D=0
M1297 405 74 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=38890 $D=0
M1298 167 75 406 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=34260 $D=0
M1299 168 75 407 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=38890 $D=0
M1300 408 76 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=34260 $D=0
M1301 409 76 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=38890 $D=0
M1302 410 406 210 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=34260 $D=0
M1303 411 407 211 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=38890 $D=0
M1304 167 410 723 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=34260 $D=0
M1305 168 411 724 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=38890 $D=0
M1306 412 723 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=34260 $D=0
M1307 413 724 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=38890 $D=0
M1308 410 75 412 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=34260 $D=0
M1309 411 75 413 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=38890 $D=0
M1310 412 408 220 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=34260 $D=0
M1311 413 409 221 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=38890 $D=0
M1312 224 414 412 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=34260 $D=0
M1313 225 415 413 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=38890 $D=0
M1314 414 77 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=34260 $D=0
M1315 415 77 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=38890 $D=0
M1316 167 78 416 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=34260 $D=0
M1317 168 78 417 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=38890 $D=0
M1318 418 79 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=34260 $D=0
M1319 419 79 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=38890 $D=0
M1320 420 416 210 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=34260 $D=0
M1321 421 417 211 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=38890 $D=0
M1322 167 420 725 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=34260 $D=0
M1323 168 421 726 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=38890 $D=0
M1324 422 725 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=34260 $D=0
M1325 423 726 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=38890 $D=0
M1326 420 78 422 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=34260 $D=0
M1327 421 78 423 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=38890 $D=0
M1328 422 418 220 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=34260 $D=0
M1329 423 419 221 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=38890 $D=0
M1330 224 424 422 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=34260 $D=0
M1331 225 425 423 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=38890 $D=0
M1332 424 80 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=34260 $D=0
M1333 425 80 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=38890 $D=0
M1334 167 81 426 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=34260 $D=0
M1335 168 81 427 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=38890 $D=0
M1336 428 82 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=34260 $D=0
M1337 429 82 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=38890 $D=0
M1338 430 426 210 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=34260 $D=0
M1339 431 427 211 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=38890 $D=0
M1340 167 430 727 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=34260 $D=0
M1341 168 431 728 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=38890 $D=0
M1342 432 727 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=34260 $D=0
M1343 433 728 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=38890 $D=0
M1344 430 81 432 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=34260 $D=0
M1345 431 81 433 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=38890 $D=0
M1346 432 428 220 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=34260 $D=0
M1347 433 429 221 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=38890 $D=0
M1348 224 434 432 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=34260 $D=0
M1349 225 435 433 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=38890 $D=0
M1350 434 83 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=34260 $D=0
M1351 435 83 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=38890 $D=0
M1352 167 84 436 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=34260 $D=0
M1353 168 84 437 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=38890 $D=0
M1354 438 85 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=34260 $D=0
M1355 439 85 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=38890 $D=0
M1356 440 436 210 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=34260 $D=0
M1357 441 437 211 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=38890 $D=0
M1358 167 440 729 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=34260 $D=0
M1359 168 441 730 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=38890 $D=0
M1360 442 729 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=34260 $D=0
M1361 443 730 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=38890 $D=0
M1362 440 84 442 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=34260 $D=0
M1363 441 84 443 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=38890 $D=0
M1364 442 438 220 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=34260 $D=0
M1365 443 439 221 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=38890 $D=0
M1366 224 444 442 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=34260 $D=0
M1367 225 445 443 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=38890 $D=0
M1368 444 86 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=34260 $D=0
M1369 445 86 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=38890 $D=0
M1370 167 87 446 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=34260 $D=0
M1371 168 87 447 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=38890 $D=0
M1372 448 88 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=34260 $D=0
M1373 449 88 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=38890 $D=0
M1374 450 446 210 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=34260 $D=0
M1375 451 447 211 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=38890 $D=0
M1376 167 450 731 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=34260 $D=0
M1377 168 451 732 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=38890 $D=0
M1378 452 731 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=34260 $D=0
M1379 453 732 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=38890 $D=0
M1380 450 87 452 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=34260 $D=0
M1381 451 87 453 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=38890 $D=0
M1382 452 448 220 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=34260 $D=0
M1383 453 449 221 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=38890 $D=0
M1384 224 454 452 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=34260 $D=0
M1385 225 455 453 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=38890 $D=0
M1386 454 89 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=34260 $D=0
M1387 455 89 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=38890 $D=0
M1388 167 90 456 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=34260 $D=0
M1389 168 90 457 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=38890 $D=0
M1390 458 91 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=34260 $D=0
M1391 459 91 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=38890 $D=0
M1392 460 456 210 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=34260 $D=0
M1393 461 457 211 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=38890 $D=0
M1394 167 460 733 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=34260 $D=0
M1395 168 461 734 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=38890 $D=0
M1396 462 733 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=34260 $D=0
M1397 463 734 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=38890 $D=0
M1398 460 90 462 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=34260 $D=0
M1399 461 90 463 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=38890 $D=0
M1400 462 458 220 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=34260 $D=0
M1401 463 459 221 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=38890 $D=0
M1402 224 464 462 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=34260 $D=0
M1403 225 465 463 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=38890 $D=0
M1404 464 92 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=34260 $D=0
M1405 465 92 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=38890 $D=0
M1406 167 93 466 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=34260 $D=0
M1407 168 93 467 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=38890 $D=0
M1408 468 94 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=34260 $D=0
M1409 469 94 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=38890 $D=0
M1410 470 466 210 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=34260 $D=0
M1411 471 467 211 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=38890 $D=0
M1412 167 470 735 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=34260 $D=0
M1413 168 471 736 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=38890 $D=0
M1414 472 735 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=34260 $D=0
M1415 473 736 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=38890 $D=0
M1416 470 93 472 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=34260 $D=0
M1417 471 93 473 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=38890 $D=0
M1418 472 468 220 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=34260 $D=0
M1419 473 469 221 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=38890 $D=0
M1420 224 474 472 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=34260 $D=0
M1421 225 475 473 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=38890 $D=0
M1422 474 95 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=34260 $D=0
M1423 475 95 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=38890 $D=0
M1424 167 96 476 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=34260 $D=0
M1425 168 96 477 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=38890 $D=0
M1426 478 97 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=34260 $D=0
M1427 479 97 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=38890 $D=0
M1428 480 476 210 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=34260 $D=0
M1429 481 477 211 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=38890 $D=0
M1430 167 480 737 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=34260 $D=0
M1431 168 481 738 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=38890 $D=0
M1432 482 737 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=34260 $D=0
M1433 483 738 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=38890 $D=0
M1434 480 96 482 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=34260 $D=0
M1435 481 96 483 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=38890 $D=0
M1436 482 478 220 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=34260 $D=0
M1437 483 479 221 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=38890 $D=0
M1438 224 484 482 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=34260 $D=0
M1439 225 485 483 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=38890 $D=0
M1440 484 98 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=34260 $D=0
M1441 485 98 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=38890 $D=0
M1442 167 99 486 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=34260 $D=0
M1443 168 99 487 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=38890 $D=0
M1444 488 100 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=34260 $D=0
M1445 489 100 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=38890 $D=0
M1446 490 486 210 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=34260 $D=0
M1447 491 487 211 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=38890 $D=0
M1448 167 490 739 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=34260 $D=0
M1449 168 491 740 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=38890 $D=0
M1450 492 739 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=34260 $D=0
M1451 493 740 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=38890 $D=0
M1452 490 99 492 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=34260 $D=0
M1453 491 99 493 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=38890 $D=0
M1454 492 488 220 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=34260 $D=0
M1455 493 489 221 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=38890 $D=0
M1456 224 494 492 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=34260 $D=0
M1457 225 495 493 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=38890 $D=0
M1458 494 101 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=34260 $D=0
M1459 495 101 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=38890 $D=0
M1460 167 102 496 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=34260 $D=0
M1461 168 102 497 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=38890 $D=0
M1462 498 103 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=34260 $D=0
M1463 499 103 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=38890 $D=0
M1464 500 496 210 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=34260 $D=0
M1465 501 497 211 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=38890 $D=0
M1466 167 500 741 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=34260 $D=0
M1467 168 501 742 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=38890 $D=0
M1468 502 741 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=34260 $D=0
M1469 503 742 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=38890 $D=0
M1470 500 102 502 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=34260 $D=0
M1471 501 102 503 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=38890 $D=0
M1472 502 498 220 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=34260 $D=0
M1473 503 499 221 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=38890 $D=0
M1474 224 504 502 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=34260 $D=0
M1475 225 505 503 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=38890 $D=0
M1476 504 104 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=34260 $D=0
M1477 505 104 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=38890 $D=0
M1478 167 105 506 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=34260 $D=0
M1479 168 105 507 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=38890 $D=0
M1480 508 106 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=34260 $D=0
M1481 509 106 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=38890 $D=0
M1482 510 506 210 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=34260 $D=0
M1483 511 507 211 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=38890 $D=0
M1484 167 510 743 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=34260 $D=0
M1485 168 511 744 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=38890 $D=0
M1486 512 743 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=34260 $D=0
M1487 513 744 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=38890 $D=0
M1488 510 105 512 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=34260 $D=0
M1489 511 105 513 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=38890 $D=0
M1490 512 508 220 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=34260 $D=0
M1491 513 509 221 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=38890 $D=0
M1492 224 514 512 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=34260 $D=0
M1493 225 515 513 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=38890 $D=0
M1494 514 107 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=34260 $D=0
M1495 515 107 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=38890 $D=0
M1496 167 108 516 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=34260 $D=0
M1497 168 108 517 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=38890 $D=0
M1498 518 109 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=34260 $D=0
M1499 519 109 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=38890 $D=0
M1500 520 516 210 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=34260 $D=0
M1501 521 517 211 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=38890 $D=0
M1502 167 520 745 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=34260 $D=0
M1503 168 521 746 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=38890 $D=0
M1504 522 745 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=34260 $D=0
M1505 523 746 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=38890 $D=0
M1506 520 108 522 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=34260 $D=0
M1507 521 108 523 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=38890 $D=0
M1508 522 518 220 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=34260 $D=0
M1509 523 519 221 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=38890 $D=0
M1510 224 524 522 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=34260 $D=0
M1511 225 525 523 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=38890 $D=0
M1512 524 110 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=34260 $D=0
M1513 525 110 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=38890 $D=0
M1514 167 111 526 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=34260 $D=0
M1515 168 111 527 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=38890 $D=0
M1516 528 112 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=34260 $D=0
M1517 529 112 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=38890 $D=0
M1518 6 528 220 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=34260 $D=0
M1519 7 529 221 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=38890 $D=0
M1520 224 526 6 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=34260 $D=0
M1521 225 527 7 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=38890 $D=0
M1522 167 532 530 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=34260 $D=0
M1523 168 533 531 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=38890 $D=0
M1524 532 113 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=34260 $D=0
M1525 533 113 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=38890 $D=0
M1526 747 220 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=34260 $D=0
M1527 748 221 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=38890 $D=0
M1528 534 532 747 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=34260 $D=0
M1529 535 533 748 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=38890 $D=0
M1530 167 534 536 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=34260 $D=0
M1531 168 535 537 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=38890 $D=0
M1532 749 536 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=34260 $D=0
M1533 750 537 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=38890 $D=0
M1534 534 530 749 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=34260 $D=0
M1535 535 531 750 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=38890 $D=0
M1536 167 540 538 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=34260 $D=0
M1537 168 541 539 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=38890 $D=0
M1538 540 113 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=34260 $D=0
M1539 541 113 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=38890 $D=0
M1540 751 224 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=34260 $D=0
M1541 752 225 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=38890 $D=0
M1542 542 540 751 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=34260 $D=0
M1543 543 541 752 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=38890 $D=0
M1544 167 542 114 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=34260 $D=0
M1545 168 543 115 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=38890 $D=0
M1546 753 114 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=34260 $D=0
M1547 754 115 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=38890 $D=0
M1548 542 538 753 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=34260 $D=0
M1549 543 539 754 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=38890 $D=0
M1550 544 116 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=34260 $D=0
M1551 545 116 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=38890 $D=0
M1552 546 116 536 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=34260 $D=0
M1553 547 116 537 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=38890 $D=0
M1554 117 544 546 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=34260 $D=0
M1555 118 545 547 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=38890 $D=0
M1556 548 119 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=34260 $D=0
M1557 549 119 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=38890 $D=0
M1558 550 119 114 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=34260 $D=0
M1559 551 119 115 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=38890 $D=0
M1560 755 548 550 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=34260 $D=0
M1561 756 549 551 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=38890 $D=0
M1562 167 114 755 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=34260 $D=0
M1563 168 115 756 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=38890 $D=0
M1564 552 120 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=34260 $D=0
M1565 553 120 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=38890 $D=0
M1566 554 120 550 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=34260 $D=0
M1567 555 120 551 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=38890 $D=0
M1568 12 552 554 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=34260 $D=0
M1569 13 553 555 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=38890 $D=0
M1570 557 556 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=34260 $D=0
M1571 558 121 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=38890 $D=0
M1572 167 561 559 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=34260 $D=0
M1573 168 562 560 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=38890 $D=0
M1574 563 546 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=34260 $D=0
M1575 564 547 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=38890 $D=0
M1576 561 546 556 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=34260 $D=0
M1577 562 547 121 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=38890 $D=0
M1578 557 563 561 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=34260 $D=0
M1579 558 564 562 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=38890 $D=0
M1580 565 559 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=34260 $D=0
M1581 566 560 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=38890 $D=0
M1582 122 559 554 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=34260 $D=0
M1583 556 560 555 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=38890 $D=0
M1584 546 565 122 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=34260 $D=0
M1585 547 566 556 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=38890 $D=0
M1586 567 122 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=34260 $D=0
M1587 568 556 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=38890 $D=0
M1588 569 559 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=34260 $D=0
M1589 570 560 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=38890 $D=0
M1590 571 559 567 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=34260 $D=0
M1591 572 560 568 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=38890 $D=0
M1592 554 569 571 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=34260 $D=0
M1593 555 570 572 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=38890 $D=0
M1594 775 546 167 167 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=33900 $D=0
M1595 776 547 168 168 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=38530 $D=0
M1596 573 554 775 167 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=33900 $D=0
M1597 574 555 776 168 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=38530 $D=0
M1598 575 571 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=34260 $D=0
M1599 576 572 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=38890 $D=0
M1600 577 546 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=34260 $D=0
M1601 578 547 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=38890 $D=0
M1602 167 554 577 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=34260 $D=0
M1603 168 555 578 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=38890 $D=0
M1604 579 546 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=34260 $D=0
M1605 580 547 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=38890 $D=0
M1606 167 554 579 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=34260 $D=0
M1607 168 555 580 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=38890 $D=0
M1608 777 546 167 167 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=34080 $D=0
M1609 778 547 168 168 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=38710 $D=0
M1610 583 554 777 167 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=34080 $D=0
M1611 584 555 778 168 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=38710 $D=0
M1612 167 579 583 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=34260 $D=0
M1613 168 580 584 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=38890 $D=0
M1614 585 127 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=34260 $D=0
M1615 586 127 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=38890 $D=0
M1616 587 127 573 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=34260 $D=0
M1617 588 127 574 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=38890 $D=0
M1618 577 585 587 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=34260 $D=0
M1619 578 586 588 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=38890 $D=0
M1620 589 127 575 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=34260 $D=0
M1621 590 127 576 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=38890 $D=0
M1622 583 585 589 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=34260 $D=0
M1623 584 586 590 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=38890 $D=0
M1624 591 128 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=34260 $D=0
M1625 592 128 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=38890 $D=0
M1626 593 128 589 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=34260 $D=0
M1627 594 128 590 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=38890 $D=0
M1628 587 591 593 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=34260 $D=0
M1629 588 592 594 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=38890 $D=0
M1630 14 593 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=34260 $D=0
M1631 15 594 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=38890 $D=0
M1632 595 129 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=34260 $D=0
M1633 596 129 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=38890 $D=0
M1634 597 129 130 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=34260 $D=0
M1635 598 129 131 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=38890 $D=0
M1636 132 595 597 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=34260 $D=0
M1637 133 596 598 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=38890 $D=0
M1638 599 129 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=34260 $D=0
M1639 600 129 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=38890 $D=0
M1640 602 129 134 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=34260 $D=0
M1641 603 129 136 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=38890 $D=0
M1642 137 599 602 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=34260 $D=0
M1643 135 600 603 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=38890 $D=0
M1644 604 129 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=34260 $D=0
M1645 605 129 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=38890 $D=0
M1646 606 129 123 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=34260 $D=0
M1647 607 129 126 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=38890 $D=0
M1648 138 604 606 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=34260 $D=0
M1649 139 605 607 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=38890 $D=0
M1650 608 129 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=34260 $D=0
M1651 609 129 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=38890 $D=0
M1652 610 129 140 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=34260 $D=0
M1653 611 129 141 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=38890 $D=0
M1654 142 608 610 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=34260 $D=0
M1655 143 609 611 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=38890 $D=0
M1656 612 129 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=34260 $D=0
M1657 613 129 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=38890 $D=0
M1658 614 129 144 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=34260 $D=0
M1659 615 129 145 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=38890 $D=0
M1660 142 612 614 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=34260 $D=0
M1661 142 613 615 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=38890 $D=0
M1662 167 546 765 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=34260 $D=0
M1663 168 547 766 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=38890 $D=0
M1664 133 765 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=34260 $D=0
M1665 130 766 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=38890 $D=0
M1666 616 146 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=34260 $D=0
M1667 617 146 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=38890 $D=0
M1668 147 146 133 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=34260 $D=0
M1669 148 146 130 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=38890 $D=0
M1670 597 616 147 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=34260 $D=0
M1671 598 617 148 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=38890 $D=0
M1672 618 149 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=34260 $D=0
M1673 619 149 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=38890 $D=0
M1674 150 149 147 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=34260 $D=0
M1675 125 149 148 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=38890 $D=0
M1676 602 618 150 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=34260 $D=0
M1677 603 619 125 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=38890 $D=0
M1678 620 151 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=34260 $D=0
M1679 621 151 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=38890 $D=0
M1680 152 151 150 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=34260 $D=0
M1681 153 151 125 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=38890 $D=0
M1682 606 620 152 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=34260 $D=0
M1683 607 621 153 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=38890 $D=0
M1684 622 154 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=34260 $D=0
M1685 623 154 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=38890 $D=0
M1686 155 154 152 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=34260 $D=0
M1687 156 154 153 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=38890 $D=0
M1688 610 622 155 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=34260 $D=0
M1689 611 623 156 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=38890 $D=0
M1690 624 157 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=34260 $D=0
M1691 625 157 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=38890 $D=0
M1692 196 157 155 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=34260 $D=0
M1693 197 157 156 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=38890 $D=0
M1694 614 624 196 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=34260 $D=0
M1695 615 625 197 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=38890 $D=0
M1696 626 158 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=34260 $D=0
M1697 627 158 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=38890 $D=0
M1698 628 158 114 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=34260 $D=0
M1699 629 158 115 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=38890 $D=0
M1700 12 626 628 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=34260 $D=0
M1701 13 627 629 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=38890 $D=0
M1702 630 536 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=34260 $D=0
M1703 631 537 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=38890 $D=0
M1704 167 628 630 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=34260 $D=0
M1705 168 629 631 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=38890 $D=0
M1706 779 536 167 167 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=34080 $D=0
M1707 780 537 168 168 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=38710 $D=0
M1708 634 628 779 167 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=34080 $D=0
M1709 635 629 780 168 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=38710 $D=0
M1710 167 630 634 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=34260 $D=0
M1711 168 631 635 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=38890 $D=0
M1712 767 159 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=34260 $D=0
M1713 768 636 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=38890 $D=0
M1714 167 634 767 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=34260 $D=0
M1715 168 635 768 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=38890 $D=0
M1716 636 767 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=34260 $D=0
M1717 160 768 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=38890 $D=0
M1718 781 536 167 167 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=33900 $D=0
M1719 782 537 168 168 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=38530 $D=0
M1720 637 639 781 167 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=33900 $D=0
M1721 638 640 782 168 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=38530 $D=0
M1722 639 628 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=34260 $D=0
M1723 640 629 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=38890 $D=0
M1724 641 637 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=34260 $D=0
M1725 642 638 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=38890 $D=0
M1726 167 159 641 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=34260 $D=0
M1727 168 636 642 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=38890 $D=0
M1728 644 161 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=34260 $D=0
M1729 645 643 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=38890 $D=0
M1730 643 641 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=34260 $D=0
M1731 162 642 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=38890 $D=0
M1732 167 644 643 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=34260 $D=0
M1733 168 645 162 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=38890 $D=0
M1734 647 646 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=34260 $D=0
M1735 648 163 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=38890 $D=0
M1736 167 651 649 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=34260 $D=0
M1737 168 652 650 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=38890 $D=0
M1738 653 117 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=34260 $D=0
M1739 654 118 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=38890 $D=0
M1740 651 117 646 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=34260 $D=0
M1741 652 118 163 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=38890 $D=0
M1742 647 653 651 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=34260 $D=0
M1743 648 654 652 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=38890 $D=0
M1744 655 649 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=34260 $D=0
M1745 656 650 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=38890 $D=0
M1746 164 649 6 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=34260 $D=0
M1747 646 650 7 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=38890 $D=0
M1748 117 655 164 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=34260 $D=0
M1749 118 656 646 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=38890 $D=0
M1750 657 164 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=34260 $D=0
M1751 658 646 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=38890 $D=0
M1752 659 649 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=34260 $D=0
M1753 660 650 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=38890 $D=0
M1754 198 649 657 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=34260 $D=0
M1755 199 650 658 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=38890 $D=0
M1756 6 659 198 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=34260 $D=0
M1757 7 660 199 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=38890 $D=0
M1758 661 165 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=34260 $D=0
M1759 662 165 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=38890 $D=0
M1760 663 165 198 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=34260 $D=0
M1761 664 165 199 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=38890 $D=0
M1762 14 661 663 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=34260 $D=0
M1763 15 662 664 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=38890 $D=0
M1764 665 166 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=34260 $D=0
M1765 666 166 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=38890 $D=0
M1766 166 166 663 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=34260 $D=0
M1767 166 166 664 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=38890 $D=0
M1768 6 665 166 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=34260 $D=0
M1769 7 666 166 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=38890 $D=0
M1770 667 113 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=34260 $D=0
M1771 668 113 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=38890 $D=0
M1772 167 667 669 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=34260 $D=0
M1773 168 668 670 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=38890 $D=0
M1774 671 113 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=34260 $D=0
M1775 672 113 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=38890 $D=0
M1776 673 669 166 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=34260 $D=0
M1777 674 670 166 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=38890 $D=0
M1778 167 673 769 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=34260 $D=0
M1779 168 674 770 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=38890 $D=0
M1780 675 769 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=34260 $D=0
M1781 676 770 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=38890 $D=0
M1782 673 667 675 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=34260 $D=0
M1783 674 668 676 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=38890 $D=0
M1784 677 671 675 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=34260 $D=0
M1785 678 672 676 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=38890 $D=0
M1786 167 681 679 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=34260 $D=0
M1787 168 682 680 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=38890 $D=0
M1788 681 113 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=34260 $D=0
M1789 682 113 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=38890 $D=0
M1790 771 677 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=34260 $D=0
M1791 772 678 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=38890 $D=0
M1792 683 681 771 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=34260 $D=0
M1793 684 682 772 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=38890 $D=0
M1794 167 683 117 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=34260 $D=0
M1795 168 684 118 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=38890 $D=0
M1796 773 117 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=34260 $D=0
M1797 774 118 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=38890 $D=0
M1798 683 679 773 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=34260 $D=0
M1799 684 680 774 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=38890 $D=0
.ENDS
***************************************
.SUBCKT ICV_39 1 2 3 4 5 6 7 9 10 11 12 13 14 15 16 17 18 19 20 21
+ 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41
+ 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61
+ 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81
+ 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101
+ 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121
+ 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141 142
+ 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162
+ 163 164 165
** N=793 EP=163 IP=1514 FDC=1800
M0 169 1 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=23750 $D=1
M1 170 1 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=28380 $D=1
M2 171 169 2 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=23750 $D=1
M3 172 170 3 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=28380 $D=1
M4 6 1 171 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=23750 $D=1
M5 7 1 172 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=28380 $D=1
M6 173 169 4 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=23750 $D=1
M7 174 170 4 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=28380 $D=1
M8 5 1 173 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=23750 $D=1
M9 5 1 174 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=28380 $D=1
M10 175 169 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=23750 $D=1
M11 176 170 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=28380 $D=1
M12 6 1 175 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=23750 $D=1
M13 7 1 176 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=28380 $D=1
M14 179 177 175 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=23750 $D=1
M15 180 178 176 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=28380 $D=1
M16 177 9 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=23750 $D=1
M17 178 9 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=28380 $D=1
M18 181 177 173 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=23750 $D=1
M19 182 178 174 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=28380 $D=1
M20 171 9 181 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=23750 $D=1
M21 172 9 182 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=28380 $D=1
M22 183 10 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=23750 $D=1
M23 184 10 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=28380 $D=1
M24 185 183 181 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=23750 $D=1
M25 186 184 182 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=28380 $D=1
M26 179 10 185 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=23750 $D=1
M27 180 10 186 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=28380 $D=1
M28 187 11 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=23750 $D=1
M29 188 11 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=28380 $D=1
M30 189 187 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=23750 $D=1
M31 190 188 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=28380 $D=1
M32 12 11 189 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=23750 $D=1
M33 13 11 190 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=28380 $D=1
M34 191 187 14 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=23750 $D=1
M35 192 188 15 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=28380 $D=1
M36 193 11 191 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=23750 $D=1
M37 194 11 192 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=28380 $D=1
M38 197 187 195 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=23750 $D=1
M39 198 188 196 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=28380 $D=1
M40 185 11 197 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=23750 $D=1
M41 186 11 198 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=28380 $D=1
M42 201 199 197 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=23750 $D=1
M43 202 200 198 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=28380 $D=1
M44 199 16 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=23750 $D=1
M45 200 16 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=28380 $D=1
M46 203 199 191 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=23750 $D=1
M47 204 200 192 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=28380 $D=1
M48 189 16 203 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=23750 $D=1
M49 190 16 204 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=28380 $D=1
M50 205 17 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=23750 $D=1
M51 206 17 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=28380 $D=1
M52 207 205 203 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=23750 $D=1
M53 208 206 204 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=28380 $D=1
M54 201 17 207 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=23750 $D=1
M55 202 17 208 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=28380 $D=1
M56 6 18 209 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=23750 $D=1
M57 7 18 210 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=28380 $D=1
M58 211 19 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=23750 $D=1
M59 212 19 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=28380 $D=1
M60 213 18 207 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=23750 $D=1
M61 214 18 208 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=28380 $D=1
M62 6 213 684 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=23750 $D=1
M63 7 214 685 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=28380 $D=1
M64 215 684 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=23750 $D=1
M65 216 685 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=28380 $D=1
M66 213 209 215 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=23750 $D=1
M67 214 210 216 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=28380 $D=1
M68 215 19 217 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=23750 $D=1
M69 216 19 218 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=28380 $D=1
M70 221 20 215 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=23750 $D=1
M71 222 20 216 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=28380 $D=1
M72 219 20 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=23750 $D=1
M73 220 20 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=28380 $D=1
M74 6 21 223 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=23750 $D=1
M75 7 21 224 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=28380 $D=1
M76 225 22 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=23750 $D=1
M77 226 22 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=28380 $D=1
M78 227 21 207 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=23750 $D=1
M79 228 21 208 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=28380 $D=1
M80 6 227 686 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=23750 $D=1
M81 7 228 687 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=28380 $D=1
M82 229 686 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=23750 $D=1
M83 230 687 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=28380 $D=1
M84 227 223 229 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=23750 $D=1
M85 228 224 230 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=28380 $D=1
M86 229 22 217 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=23750 $D=1
M87 230 22 218 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=28380 $D=1
M88 221 23 229 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=23750 $D=1
M89 222 23 230 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=28380 $D=1
M90 231 23 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=23750 $D=1
M91 232 23 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=28380 $D=1
M92 6 24 233 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=23750 $D=1
M93 7 24 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=28380 $D=1
M94 235 25 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=23750 $D=1
M95 236 25 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=28380 $D=1
M96 237 24 207 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=23750 $D=1
M97 238 24 208 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=28380 $D=1
M98 6 237 688 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=23750 $D=1
M99 7 238 689 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=28380 $D=1
M100 239 688 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=23750 $D=1
M101 240 689 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=28380 $D=1
M102 237 233 239 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=23750 $D=1
M103 238 234 240 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=28380 $D=1
M104 239 25 217 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=23750 $D=1
M105 240 25 218 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=28380 $D=1
M106 221 26 239 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=23750 $D=1
M107 222 26 240 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=28380 $D=1
M108 241 26 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=23750 $D=1
M109 242 26 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=28380 $D=1
M110 6 27 243 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=23750 $D=1
M111 7 27 244 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=28380 $D=1
M112 245 28 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=23750 $D=1
M113 246 28 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=28380 $D=1
M114 247 27 207 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=23750 $D=1
M115 248 27 208 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=28380 $D=1
M116 6 247 690 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=23750 $D=1
M117 7 248 691 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=28380 $D=1
M118 249 690 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=23750 $D=1
M119 250 691 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=28380 $D=1
M120 247 243 249 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=23750 $D=1
M121 248 244 250 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=28380 $D=1
M122 249 28 217 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=23750 $D=1
M123 250 28 218 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=28380 $D=1
M124 221 29 249 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=23750 $D=1
M125 222 29 250 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=28380 $D=1
M126 251 29 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=23750 $D=1
M127 252 29 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=28380 $D=1
M128 6 30 253 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=23750 $D=1
M129 7 30 254 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=28380 $D=1
M130 255 31 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=23750 $D=1
M131 256 31 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=28380 $D=1
M132 257 30 207 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=23750 $D=1
M133 258 30 208 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=28380 $D=1
M134 6 257 692 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=23750 $D=1
M135 7 258 693 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=28380 $D=1
M136 259 692 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=23750 $D=1
M137 260 693 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=28380 $D=1
M138 257 253 259 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=23750 $D=1
M139 258 254 260 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=28380 $D=1
M140 259 31 217 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=23750 $D=1
M141 260 31 218 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=28380 $D=1
M142 221 32 259 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=23750 $D=1
M143 222 32 260 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=28380 $D=1
M144 261 32 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=23750 $D=1
M145 262 32 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=28380 $D=1
M146 6 33 263 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=23750 $D=1
M147 7 33 264 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=28380 $D=1
M148 265 34 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=23750 $D=1
M149 266 34 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=28380 $D=1
M150 267 33 207 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=23750 $D=1
M151 268 33 208 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=28380 $D=1
M152 6 267 694 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=23750 $D=1
M153 7 268 695 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=28380 $D=1
M154 269 694 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=23750 $D=1
M155 270 695 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=28380 $D=1
M156 267 263 269 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=23750 $D=1
M157 268 264 270 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=28380 $D=1
M158 269 34 217 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=23750 $D=1
M159 270 34 218 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=28380 $D=1
M160 221 35 269 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=23750 $D=1
M161 222 35 270 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=28380 $D=1
M162 271 35 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=23750 $D=1
M163 272 35 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=28380 $D=1
M164 6 36 273 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=23750 $D=1
M165 7 36 274 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=28380 $D=1
M166 275 37 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=23750 $D=1
M167 276 37 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=28380 $D=1
M168 277 36 207 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=23750 $D=1
M169 278 36 208 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=28380 $D=1
M170 6 277 696 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=23750 $D=1
M171 7 278 697 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=28380 $D=1
M172 279 696 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=23750 $D=1
M173 280 697 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=28380 $D=1
M174 277 273 279 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=23750 $D=1
M175 278 274 280 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=28380 $D=1
M176 279 37 217 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=23750 $D=1
M177 280 37 218 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=28380 $D=1
M178 221 38 279 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=23750 $D=1
M179 222 38 280 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=28380 $D=1
M180 281 38 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=23750 $D=1
M181 282 38 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=28380 $D=1
M182 6 39 283 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=23750 $D=1
M183 7 39 284 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=28380 $D=1
M184 285 40 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=23750 $D=1
M185 286 40 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=28380 $D=1
M186 287 39 207 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=23750 $D=1
M187 288 39 208 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=28380 $D=1
M188 6 287 698 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=23750 $D=1
M189 7 288 699 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=28380 $D=1
M190 289 698 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=23750 $D=1
M191 290 699 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=28380 $D=1
M192 287 283 289 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=23750 $D=1
M193 288 284 290 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=28380 $D=1
M194 289 40 217 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=23750 $D=1
M195 290 40 218 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=28380 $D=1
M196 221 41 289 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=23750 $D=1
M197 222 41 290 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=28380 $D=1
M198 291 41 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=23750 $D=1
M199 292 41 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=28380 $D=1
M200 6 42 293 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=23750 $D=1
M201 7 42 294 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=28380 $D=1
M202 295 43 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=23750 $D=1
M203 296 43 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=28380 $D=1
M204 297 42 207 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=23750 $D=1
M205 298 42 208 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=28380 $D=1
M206 6 297 700 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=23750 $D=1
M207 7 298 701 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=28380 $D=1
M208 299 700 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=23750 $D=1
M209 300 701 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=28380 $D=1
M210 297 293 299 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=23750 $D=1
M211 298 294 300 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=28380 $D=1
M212 299 43 217 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=23750 $D=1
M213 300 43 218 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=28380 $D=1
M214 221 44 299 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=23750 $D=1
M215 222 44 300 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=28380 $D=1
M216 301 44 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=23750 $D=1
M217 302 44 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=28380 $D=1
M218 6 45 303 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=23750 $D=1
M219 7 45 304 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=28380 $D=1
M220 305 46 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=23750 $D=1
M221 306 46 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=28380 $D=1
M222 307 45 207 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=23750 $D=1
M223 308 45 208 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=28380 $D=1
M224 6 307 702 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=23750 $D=1
M225 7 308 703 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=28380 $D=1
M226 309 702 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=23750 $D=1
M227 310 703 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=28380 $D=1
M228 307 303 309 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=23750 $D=1
M229 308 304 310 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=28380 $D=1
M230 309 46 217 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=23750 $D=1
M231 310 46 218 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=28380 $D=1
M232 221 47 309 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=23750 $D=1
M233 222 47 310 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=28380 $D=1
M234 311 47 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=23750 $D=1
M235 312 47 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=28380 $D=1
M236 6 48 313 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=23750 $D=1
M237 7 48 314 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=28380 $D=1
M238 315 49 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=23750 $D=1
M239 316 49 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=28380 $D=1
M240 317 48 207 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=23750 $D=1
M241 318 48 208 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=28380 $D=1
M242 6 317 704 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=23750 $D=1
M243 7 318 705 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=28380 $D=1
M244 319 704 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=23750 $D=1
M245 320 705 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=28380 $D=1
M246 317 313 319 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=23750 $D=1
M247 318 314 320 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=28380 $D=1
M248 319 49 217 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=23750 $D=1
M249 320 49 218 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=28380 $D=1
M250 221 50 319 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=23750 $D=1
M251 222 50 320 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=28380 $D=1
M252 321 50 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=23750 $D=1
M253 322 50 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=28380 $D=1
M254 6 51 323 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=23750 $D=1
M255 7 51 324 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=28380 $D=1
M256 325 52 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=23750 $D=1
M257 326 52 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=28380 $D=1
M258 327 51 207 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=23750 $D=1
M259 328 51 208 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=28380 $D=1
M260 6 327 706 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=23750 $D=1
M261 7 328 707 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=28380 $D=1
M262 329 706 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=23750 $D=1
M263 330 707 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=28380 $D=1
M264 327 323 329 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=23750 $D=1
M265 328 324 330 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=28380 $D=1
M266 329 52 217 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=23750 $D=1
M267 330 52 218 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=28380 $D=1
M268 221 53 329 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=23750 $D=1
M269 222 53 330 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=28380 $D=1
M270 331 53 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=23750 $D=1
M271 332 53 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=28380 $D=1
M272 6 54 333 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=23750 $D=1
M273 7 54 334 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=28380 $D=1
M274 335 55 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=23750 $D=1
M275 336 55 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=28380 $D=1
M276 337 54 207 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=23750 $D=1
M277 338 54 208 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=28380 $D=1
M278 6 337 708 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=23750 $D=1
M279 7 338 709 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=28380 $D=1
M280 339 708 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=23750 $D=1
M281 340 709 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=28380 $D=1
M282 337 333 339 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=23750 $D=1
M283 338 334 340 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=28380 $D=1
M284 339 55 217 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=23750 $D=1
M285 340 55 218 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=28380 $D=1
M286 221 56 339 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=23750 $D=1
M287 222 56 340 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=28380 $D=1
M288 341 56 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=23750 $D=1
M289 342 56 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=28380 $D=1
M290 6 57 343 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=23750 $D=1
M291 7 57 344 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=28380 $D=1
M292 345 58 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=23750 $D=1
M293 346 58 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=28380 $D=1
M294 347 57 207 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=23750 $D=1
M295 348 57 208 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=28380 $D=1
M296 6 347 710 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=23750 $D=1
M297 7 348 711 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=28380 $D=1
M298 349 710 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=23750 $D=1
M299 350 711 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=28380 $D=1
M300 347 343 349 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=23750 $D=1
M301 348 344 350 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=28380 $D=1
M302 349 58 217 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=23750 $D=1
M303 350 58 218 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=28380 $D=1
M304 221 59 349 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=23750 $D=1
M305 222 59 350 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=28380 $D=1
M306 351 59 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=23750 $D=1
M307 352 59 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=28380 $D=1
M308 6 60 353 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=23750 $D=1
M309 7 60 354 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=28380 $D=1
M310 355 61 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=23750 $D=1
M311 356 61 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=28380 $D=1
M312 357 60 207 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=23750 $D=1
M313 358 60 208 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=28380 $D=1
M314 6 357 712 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=23750 $D=1
M315 7 358 713 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=28380 $D=1
M316 359 712 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=23750 $D=1
M317 360 713 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=28380 $D=1
M318 357 353 359 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=23750 $D=1
M319 358 354 360 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=28380 $D=1
M320 359 61 217 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=23750 $D=1
M321 360 61 218 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=28380 $D=1
M322 221 62 359 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=23750 $D=1
M323 222 62 360 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=28380 $D=1
M324 361 62 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=23750 $D=1
M325 362 62 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=28380 $D=1
M326 6 63 363 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=23750 $D=1
M327 7 63 364 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=28380 $D=1
M328 365 64 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=23750 $D=1
M329 366 64 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=28380 $D=1
M330 367 63 207 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=23750 $D=1
M331 368 63 208 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=28380 $D=1
M332 6 367 714 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=23750 $D=1
M333 7 368 715 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=28380 $D=1
M334 369 714 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=23750 $D=1
M335 370 715 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=28380 $D=1
M336 367 363 369 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=23750 $D=1
M337 368 364 370 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=28380 $D=1
M338 369 64 217 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=23750 $D=1
M339 370 64 218 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=28380 $D=1
M340 221 65 369 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=23750 $D=1
M341 222 65 370 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=28380 $D=1
M342 371 65 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=23750 $D=1
M343 372 65 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=28380 $D=1
M344 6 66 373 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=23750 $D=1
M345 7 66 374 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=28380 $D=1
M346 375 67 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=23750 $D=1
M347 376 67 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=28380 $D=1
M348 377 66 207 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=23750 $D=1
M349 378 66 208 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=28380 $D=1
M350 6 377 716 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=23750 $D=1
M351 7 378 717 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=28380 $D=1
M352 379 716 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=23750 $D=1
M353 380 717 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=28380 $D=1
M354 377 373 379 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=23750 $D=1
M355 378 374 380 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=28380 $D=1
M356 379 67 217 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=23750 $D=1
M357 380 67 218 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=28380 $D=1
M358 221 68 379 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=23750 $D=1
M359 222 68 380 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=28380 $D=1
M360 381 68 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=23750 $D=1
M361 382 68 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=28380 $D=1
M362 6 69 383 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=23750 $D=1
M363 7 69 384 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=28380 $D=1
M364 385 70 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=23750 $D=1
M365 386 70 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=28380 $D=1
M366 387 69 207 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=23750 $D=1
M367 388 69 208 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=28380 $D=1
M368 6 387 718 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=23750 $D=1
M369 7 388 719 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=28380 $D=1
M370 389 718 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=23750 $D=1
M371 390 719 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=28380 $D=1
M372 387 383 389 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=23750 $D=1
M373 388 384 390 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=28380 $D=1
M374 389 70 217 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=23750 $D=1
M375 390 70 218 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=28380 $D=1
M376 221 71 389 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=23750 $D=1
M377 222 71 390 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=28380 $D=1
M378 391 71 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=23750 $D=1
M379 392 71 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=28380 $D=1
M380 6 72 393 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=23750 $D=1
M381 7 72 394 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=28380 $D=1
M382 395 73 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=23750 $D=1
M383 396 73 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=28380 $D=1
M384 397 72 207 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=23750 $D=1
M385 398 72 208 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=28380 $D=1
M386 6 397 720 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=23750 $D=1
M387 7 398 721 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=28380 $D=1
M388 399 720 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=23750 $D=1
M389 400 721 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=28380 $D=1
M390 397 393 399 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=23750 $D=1
M391 398 394 400 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=28380 $D=1
M392 399 73 217 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=23750 $D=1
M393 400 73 218 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=28380 $D=1
M394 221 74 399 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=23750 $D=1
M395 222 74 400 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=28380 $D=1
M396 401 74 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=23750 $D=1
M397 402 74 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=28380 $D=1
M398 6 75 403 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=23750 $D=1
M399 7 75 404 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=28380 $D=1
M400 405 76 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=23750 $D=1
M401 406 76 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=28380 $D=1
M402 407 75 207 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=23750 $D=1
M403 408 75 208 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=28380 $D=1
M404 6 407 722 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=23750 $D=1
M405 7 408 723 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=28380 $D=1
M406 409 722 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=23750 $D=1
M407 410 723 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=28380 $D=1
M408 407 403 409 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=23750 $D=1
M409 408 404 410 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=28380 $D=1
M410 409 76 217 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=23750 $D=1
M411 410 76 218 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=28380 $D=1
M412 221 77 409 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=23750 $D=1
M413 222 77 410 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=28380 $D=1
M414 411 77 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=23750 $D=1
M415 412 77 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=28380 $D=1
M416 6 78 413 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=23750 $D=1
M417 7 78 414 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=28380 $D=1
M418 415 79 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=23750 $D=1
M419 416 79 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=28380 $D=1
M420 417 78 207 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=23750 $D=1
M421 418 78 208 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=28380 $D=1
M422 6 417 724 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=23750 $D=1
M423 7 418 725 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=28380 $D=1
M424 419 724 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=23750 $D=1
M425 420 725 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=28380 $D=1
M426 417 413 419 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=23750 $D=1
M427 418 414 420 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=28380 $D=1
M428 419 79 217 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=23750 $D=1
M429 420 79 218 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=28380 $D=1
M430 221 80 419 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=23750 $D=1
M431 222 80 420 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=28380 $D=1
M432 421 80 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=23750 $D=1
M433 422 80 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=28380 $D=1
M434 6 81 423 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=23750 $D=1
M435 7 81 424 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=28380 $D=1
M436 425 82 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=23750 $D=1
M437 426 82 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=28380 $D=1
M438 427 81 207 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=23750 $D=1
M439 428 81 208 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=28380 $D=1
M440 6 427 726 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=23750 $D=1
M441 7 428 727 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=28380 $D=1
M442 429 726 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=23750 $D=1
M443 430 727 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=28380 $D=1
M444 427 423 429 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=23750 $D=1
M445 428 424 430 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=28380 $D=1
M446 429 82 217 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=23750 $D=1
M447 430 82 218 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=28380 $D=1
M448 221 83 429 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=23750 $D=1
M449 222 83 430 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=28380 $D=1
M450 431 83 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=23750 $D=1
M451 432 83 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=28380 $D=1
M452 6 84 433 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=23750 $D=1
M453 7 84 434 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=28380 $D=1
M454 435 85 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=23750 $D=1
M455 436 85 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=28380 $D=1
M456 437 84 207 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=23750 $D=1
M457 438 84 208 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=28380 $D=1
M458 6 437 728 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=23750 $D=1
M459 7 438 729 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=28380 $D=1
M460 439 728 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=23750 $D=1
M461 440 729 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=28380 $D=1
M462 437 433 439 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=23750 $D=1
M463 438 434 440 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=28380 $D=1
M464 439 85 217 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=23750 $D=1
M465 440 85 218 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=28380 $D=1
M466 221 86 439 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=23750 $D=1
M467 222 86 440 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=28380 $D=1
M468 441 86 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=23750 $D=1
M469 442 86 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=28380 $D=1
M470 6 87 443 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=23750 $D=1
M471 7 87 444 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=28380 $D=1
M472 445 88 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=23750 $D=1
M473 446 88 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=28380 $D=1
M474 447 87 207 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=23750 $D=1
M475 448 87 208 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=28380 $D=1
M476 6 447 730 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=23750 $D=1
M477 7 448 731 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=28380 $D=1
M478 449 730 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=23750 $D=1
M479 450 731 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=28380 $D=1
M480 447 443 449 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=23750 $D=1
M481 448 444 450 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=28380 $D=1
M482 449 88 217 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=23750 $D=1
M483 450 88 218 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=28380 $D=1
M484 221 89 449 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=23750 $D=1
M485 222 89 450 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=28380 $D=1
M486 451 89 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=23750 $D=1
M487 452 89 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=28380 $D=1
M488 6 90 453 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=23750 $D=1
M489 7 90 454 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=28380 $D=1
M490 455 91 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=23750 $D=1
M491 456 91 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=28380 $D=1
M492 457 90 207 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=23750 $D=1
M493 458 90 208 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=28380 $D=1
M494 6 457 732 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=23750 $D=1
M495 7 458 733 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=28380 $D=1
M496 459 732 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=23750 $D=1
M497 460 733 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=28380 $D=1
M498 457 453 459 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=23750 $D=1
M499 458 454 460 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=28380 $D=1
M500 459 91 217 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=23750 $D=1
M501 460 91 218 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=28380 $D=1
M502 221 92 459 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=23750 $D=1
M503 222 92 460 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=28380 $D=1
M504 461 92 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=23750 $D=1
M505 462 92 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=28380 $D=1
M506 6 93 463 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=23750 $D=1
M507 7 93 464 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=28380 $D=1
M508 465 94 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=23750 $D=1
M509 466 94 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=28380 $D=1
M510 467 93 207 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=23750 $D=1
M511 468 93 208 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=28380 $D=1
M512 6 467 734 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=23750 $D=1
M513 7 468 735 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=28380 $D=1
M514 469 734 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=23750 $D=1
M515 470 735 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=28380 $D=1
M516 467 463 469 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=23750 $D=1
M517 468 464 470 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=28380 $D=1
M518 469 94 217 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=23750 $D=1
M519 470 94 218 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=28380 $D=1
M520 221 95 469 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=23750 $D=1
M521 222 95 470 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=28380 $D=1
M522 471 95 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=23750 $D=1
M523 472 95 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=28380 $D=1
M524 6 96 473 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=23750 $D=1
M525 7 96 474 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=28380 $D=1
M526 475 97 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=23750 $D=1
M527 476 97 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=28380 $D=1
M528 477 96 207 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=23750 $D=1
M529 478 96 208 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=28380 $D=1
M530 6 477 736 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=23750 $D=1
M531 7 478 737 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=28380 $D=1
M532 479 736 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=23750 $D=1
M533 480 737 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=28380 $D=1
M534 477 473 479 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=23750 $D=1
M535 478 474 480 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=28380 $D=1
M536 479 97 217 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=23750 $D=1
M537 480 97 218 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=28380 $D=1
M538 221 98 479 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=23750 $D=1
M539 222 98 480 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=28380 $D=1
M540 481 98 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=23750 $D=1
M541 482 98 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=28380 $D=1
M542 6 99 483 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=23750 $D=1
M543 7 99 484 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=28380 $D=1
M544 485 100 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=23750 $D=1
M545 486 100 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=28380 $D=1
M546 487 99 207 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=23750 $D=1
M547 488 99 208 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=28380 $D=1
M548 6 487 738 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=23750 $D=1
M549 7 488 739 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=28380 $D=1
M550 489 738 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=23750 $D=1
M551 490 739 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=28380 $D=1
M552 487 483 489 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=23750 $D=1
M553 488 484 490 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=28380 $D=1
M554 489 100 217 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=23750 $D=1
M555 490 100 218 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=28380 $D=1
M556 221 101 489 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=23750 $D=1
M557 222 101 490 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=28380 $D=1
M558 491 101 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=23750 $D=1
M559 492 101 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=28380 $D=1
M560 6 102 493 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=23750 $D=1
M561 7 102 494 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=28380 $D=1
M562 495 103 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=23750 $D=1
M563 496 103 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=28380 $D=1
M564 497 102 207 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=23750 $D=1
M565 498 102 208 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=28380 $D=1
M566 6 497 740 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=23750 $D=1
M567 7 498 741 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=28380 $D=1
M568 499 740 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=23750 $D=1
M569 500 741 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=28380 $D=1
M570 497 493 499 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=23750 $D=1
M571 498 494 500 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=28380 $D=1
M572 499 103 217 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=23750 $D=1
M573 500 103 218 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=28380 $D=1
M574 221 104 499 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=23750 $D=1
M575 222 104 500 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=28380 $D=1
M576 501 104 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=23750 $D=1
M577 502 104 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=28380 $D=1
M578 6 105 503 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=23750 $D=1
M579 7 105 504 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=28380 $D=1
M580 505 106 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=23750 $D=1
M581 506 106 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=28380 $D=1
M582 507 105 207 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=23750 $D=1
M583 508 105 208 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=28380 $D=1
M584 6 507 742 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=23750 $D=1
M585 7 508 743 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=28380 $D=1
M586 509 742 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=23750 $D=1
M587 510 743 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=28380 $D=1
M588 507 503 509 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=23750 $D=1
M589 508 504 510 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=28380 $D=1
M590 509 106 217 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=23750 $D=1
M591 510 106 218 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=28380 $D=1
M592 221 107 509 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=23750 $D=1
M593 222 107 510 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=28380 $D=1
M594 511 107 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=23750 $D=1
M595 512 107 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=28380 $D=1
M596 6 108 513 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=23750 $D=1
M597 7 108 514 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=28380 $D=1
M598 515 109 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=23750 $D=1
M599 516 109 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=28380 $D=1
M600 517 108 207 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=23750 $D=1
M601 518 108 208 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=28380 $D=1
M602 6 517 744 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=23750 $D=1
M603 7 518 745 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=28380 $D=1
M604 519 744 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=23750 $D=1
M605 520 745 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=28380 $D=1
M606 517 513 519 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=23750 $D=1
M607 518 514 520 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=28380 $D=1
M608 519 109 217 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=23750 $D=1
M609 520 109 218 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=28380 $D=1
M610 221 110 519 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=23750 $D=1
M611 222 110 520 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=28380 $D=1
M612 521 110 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=23750 $D=1
M613 522 110 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=28380 $D=1
M614 6 111 523 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=23750 $D=1
M615 7 111 524 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=28380 $D=1
M616 525 112 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=23750 $D=1
M617 526 112 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=28380 $D=1
M618 6 112 217 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=23750 $D=1
M619 7 112 218 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=28380 $D=1
M620 221 111 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=23750 $D=1
M621 222 111 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=28380 $D=1
M622 6 529 527 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=23750 $D=1
M623 7 530 528 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=28380 $D=1
M624 529 113 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=23750 $D=1
M625 530 113 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=28380 $D=1
M626 746 217 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=23750 $D=1
M627 747 218 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=28380 $D=1
M628 531 527 746 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=23750 $D=1
M629 532 528 747 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=28380 $D=1
M630 6 531 533 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=23750 $D=1
M631 7 532 534 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=28380 $D=1
M632 748 533 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=23750 $D=1
M633 749 534 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=28380 $D=1
M634 531 529 748 6 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=23750 $D=1
M635 532 530 749 7 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=28380 $D=1
M636 6 537 535 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=23750 $D=1
M637 7 538 536 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=28380 $D=1
M638 537 113 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=23750 $D=1
M639 538 113 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=28380 $D=1
M640 750 221 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=23750 $D=1
M641 751 222 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=28380 $D=1
M642 539 535 750 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=23750 $D=1
M643 540 536 751 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=28380 $D=1
M644 6 539 114 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=23750 $D=1
M645 7 540 115 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=28380 $D=1
M646 752 114 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=23750 $D=1
M647 753 115 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=28380 $D=1
M648 539 537 752 6 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=23750 $D=1
M649 540 538 753 7 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=28380 $D=1
M650 541 116 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=23750 $D=1
M651 542 116 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=28380 $D=1
M652 543 541 533 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=23750 $D=1
M653 544 542 534 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=28380 $D=1
M654 117 116 543 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=23750 $D=1
M655 118 116 544 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=28380 $D=1
M656 545 119 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=23750 $D=1
M657 546 119 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=28380 $D=1
M658 547 545 114 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=23750 $D=1
M659 548 546 115 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=28380 $D=1
M660 754 119 547 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=23750 $D=1
M661 755 119 548 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=28380 $D=1
M662 6 114 754 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=23750 $D=1
M663 7 115 755 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=28380 $D=1
M664 549 120 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=23750 $D=1
M665 550 120 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=28380 $D=1
M666 551 549 547 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=23750 $D=1
M667 552 550 548 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=28380 $D=1
M668 12 120 551 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=23750 $D=1
M669 13 120 552 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=28380 $D=1
M670 555 553 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=23750 $D=1
M671 556 554 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=28380 $D=1
M672 6 559 557 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=23750 $D=1
M673 7 560 558 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=28380 $D=1
M674 561 543 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=23750 $D=1
M675 562 544 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=28380 $D=1
M676 559 561 553 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=23750 $D=1
M677 560 562 554 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=28380 $D=1
M678 555 543 559 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=23750 $D=1
M679 556 544 560 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=28380 $D=1
M680 563 557 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=23750 $D=1
M681 564 558 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=28380 $D=1
M682 121 563 551 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=23750 $D=1
M683 553 564 552 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=28380 $D=1
M684 543 557 121 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=23750 $D=1
M685 544 558 553 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=28380 $D=1
M686 565 121 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=23750 $D=1
M687 566 553 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=28380 $D=1
M688 567 557 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=23750 $D=1
M689 568 558 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=28380 $D=1
M690 569 567 565 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=23750 $D=1
M691 570 568 566 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=28380 $D=1
M692 551 557 569 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=23750 $D=1
M693 552 558 570 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=28380 $D=1
M694 571 543 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=23750 $D=1
M695 572 544 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=28380 $D=1
M696 6 551 571 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=23750 $D=1
M697 7 552 572 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=28380 $D=1
M698 573 569 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=23750 $D=1
M699 574 570 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=28380 $D=1
M700 782 543 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=23750 $D=1
M701 783 544 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=28380 $D=1
M702 575 551 782 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=23750 $D=1
M703 576 552 783 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=28380 $D=1
M704 784 543 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=23750 $D=1
M705 785 544 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=28380 $D=1
M706 577 551 784 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=23750 $D=1
M707 578 552 785 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=28380 $D=1
M708 581 543 579 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=23750 $D=1
M709 582 544 580 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=28380 $D=1
M710 579 551 581 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=23750 $D=1
M711 580 552 582 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=28380 $D=1
M712 6 577 579 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=23750 $D=1
M713 7 578 580 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=28380 $D=1
M714 583 126 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=23750 $D=1
M715 584 126 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=28380 $D=1
M716 585 583 571 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=23750 $D=1
M717 586 584 572 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=28380 $D=1
M718 575 126 585 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=23750 $D=1
M719 576 126 586 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=28380 $D=1
M720 587 583 573 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=23750 $D=1
M721 588 584 574 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=28380 $D=1
M722 581 126 587 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=23750 $D=1
M723 582 126 588 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=28380 $D=1
M724 589 127 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=23750 $D=1
M725 590 127 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=28380 $D=1
M726 591 589 587 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=23750 $D=1
M727 592 590 588 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=28380 $D=1
M728 585 127 591 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=23750 $D=1
M729 586 127 592 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=28380 $D=1
M730 14 591 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=23750 $D=1
M731 15 592 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=28380 $D=1
M732 593 128 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=23750 $D=1
M733 594 128 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=28380 $D=1
M734 595 593 129 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=23750 $D=1
M735 596 594 130 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=28380 $D=1
M736 131 128 595 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=23750 $D=1
M737 132 128 596 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=28380 $D=1
M738 597 128 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=23750 $D=1
M739 598 128 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=28380 $D=1
M740 600 597 133 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=23750 $D=1
M741 601 598 135 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=28380 $D=1
M742 136 128 600 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=23750 $D=1
M743 134 128 601 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=28380 $D=1
M744 602 128 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=23750 $D=1
M745 603 128 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=28380 $D=1
M746 604 602 125 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=23750 $D=1
M747 605 603 124 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=28380 $D=1
M748 137 128 604 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=23750 $D=1
M749 138 128 605 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=28380 $D=1
M750 606 128 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=23750 $D=1
M751 607 128 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=28380 $D=1
M752 608 606 139 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=23750 $D=1
M753 609 607 140 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=28380 $D=1
M754 141 128 608 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=23750 $D=1
M755 141 128 609 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=28380 $D=1
M756 610 128 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=23750 $D=1
M757 611 128 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=28380 $D=1
M758 612 610 142 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=23750 $D=1
M759 613 611 143 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=28380 $D=1
M760 141 128 612 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=23750 $D=1
M761 141 128 613 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=28380 $D=1
M762 6 543 764 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=23750 $D=1
M763 7 544 765 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=28380 $D=1
M764 132 764 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=23750 $D=1
M765 129 765 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=28380 $D=1
M766 614 144 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=23750 $D=1
M767 615 144 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=28380 $D=1
M768 145 614 132 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=23750 $D=1
M769 146 615 129 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=28380 $D=1
M770 595 144 145 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=23750 $D=1
M771 596 144 146 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=28380 $D=1
M772 616 147 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=23750 $D=1
M773 617 147 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=28380 $D=1
M774 148 616 145 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=23750 $D=1
M775 123 617 146 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=28380 $D=1
M776 600 147 148 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=23750 $D=1
M777 601 147 123 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=28380 $D=1
M778 618 149 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=23750 $D=1
M779 619 149 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=28380 $D=1
M780 150 618 148 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=23750 $D=1
M781 151 619 123 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=28380 $D=1
M782 604 149 150 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=23750 $D=1
M783 605 149 151 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=28380 $D=1
M784 620 152 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=23750 $D=1
M785 621 152 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=28380 $D=1
M786 153 620 150 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=23750 $D=1
M787 154 621 151 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=28380 $D=1
M788 608 152 153 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=23750 $D=1
M789 609 152 154 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=28380 $D=1
M790 622 155 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=23750 $D=1
M791 623 155 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=28380 $D=1
M792 193 622 153 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=23750 $D=1
M793 194 623 154 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=28380 $D=1
M794 612 155 193 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=23750 $D=1
M795 613 155 194 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=28380 $D=1
M796 624 156 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=23750 $D=1
M797 625 156 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=28380 $D=1
M798 626 624 114 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=23750 $D=1
M799 627 625 115 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=28380 $D=1
M800 12 156 626 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=23750 $D=1
M801 13 156 627 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=28380 $D=1
M802 786 533 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=23750 $D=1
M803 787 534 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=28380 $D=1
M804 628 626 786 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=23750 $D=1
M805 629 627 787 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=28380 $D=1
M806 632 533 630 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=23750 $D=1
M807 633 534 631 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=28380 $D=1
M808 630 626 632 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=23750 $D=1
M809 631 627 633 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=28380 $D=1
M810 6 628 630 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=23750 $D=1
M811 7 629 631 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=28380 $D=1
M812 788 157 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=23750 $D=1
M813 789 634 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=28380 $D=1
M814 766 632 788 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=23750 $D=1
M815 767 633 789 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=28380 $D=1
M816 634 766 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=23750 $D=1
M817 635 767 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=28380 $D=1
M818 636 533 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=23750 $D=1
M819 637 534 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=28380 $D=1
M820 6 638 636 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=23750 $D=1
M821 7 639 637 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=28380 $D=1
M822 638 626 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=23750 $D=1
M823 639 627 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=28380 $D=1
M824 790 636 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=23750 $D=1
M825 791 637 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=28380 $D=1
M826 640 157 790 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=23750 $D=1
M827 641 634 791 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=28380 $D=1
M828 643 158 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=23750 $D=1
M829 644 642 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=28380 $D=1
M830 792 640 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=23750 $D=1
M831 793 641 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=28380 $D=1
M832 642 643 792 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=23750 $D=1
M833 159 644 793 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=28380 $D=1
M834 646 645 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=23750 $D=1
M835 647 160 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=28380 $D=1
M836 6 650 648 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=23750 $D=1
M837 7 651 649 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=28380 $D=1
M838 652 117 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=23750 $D=1
M839 653 118 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=28380 $D=1
M840 650 652 645 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=23750 $D=1
M841 651 653 160 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=28380 $D=1
M842 646 117 650 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=23750 $D=1
M843 647 118 651 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=28380 $D=1
M844 654 648 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=23750 $D=1
M845 655 649 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=28380 $D=1
M846 161 654 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=23750 $D=1
M847 645 655 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=28380 $D=1
M848 117 648 161 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=23750 $D=1
M849 118 649 645 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=28380 $D=1
M850 656 161 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=23750 $D=1
M851 657 645 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=28380 $D=1
M852 658 648 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=23750 $D=1
M853 659 649 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=28380 $D=1
M854 195 658 656 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=23750 $D=1
M855 196 659 657 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=28380 $D=1
M856 6 648 195 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=23750 $D=1
M857 7 649 196 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=28380 $D=1
M858 660 162 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=23750 $D=1
M859 661 162 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=28380 $D=1
M860 662 660 195 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=23750 $D=1
M861 663 661 196 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=28380 $D=1
M862 14 162 662 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=23750 $D=1
M863 15 162 663 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=28380 $D=1
M864 664 163 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=23750 $D=1
M865 665 163 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=28380 $D=1
M866 163 664 662 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=23750 $D=1
M867 163 665 663 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=28380 $D=1
M868 6 163 163 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=23750 $D=1
M869 7 163 163 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=28380 $D=1
M870 666 113 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=23750 $D=1
M871 667 113 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=28380 $D=1
M872 6 666 668 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=23750 $D=1
M873 7 667 669 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=28380 $D=1
M874 670 113 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=23750 $D=1
M875 671 113 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=28380 $D=1
M876 672 666 163 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=23750 $D=1
M877 673 667 163 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=28380 $D=1
M878 6 672 768 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=23750 $D=1
M879 7 673 769 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=28380 $D=1
M880 674 768 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=23750 $D=1
M881 675 769 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=28380 $D=1
M882 672 668 674 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=23750 $D=1
M883 673 669 675 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=28380 $D=1
M884 676 113 674 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=23750 $D=1
M885 677 113 675 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=28380 $D=1
M886 6 680 678 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=23750 $D=1
M887 7 681 679 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=28380 $D=1
M888 680 113 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=23750 $D=1
M889 681 113 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=28380 $D=1
M890 770 676 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=23750 $D=1
M891 771 677 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=28380 $D=1
M892 682 678 770 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=23750 $D=1
M893 683 679 771 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=28380 $D=1
M894 6 682 117 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=23750 $D=1
M895 7 683 118 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=28380 $D=1
M896 772 117 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=23750 $D=1
M897 773 118 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=28380 $D=1
M898 682 680 772 6 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=23750 $D=1
M899 683 681 773 7 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=28380 $D=1
M900 169 1 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=25000 $D=0
M901 170 1 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=29630 $D=0
M902 171 1 2 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=25000 $D=0
M903 172 1 3 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=29630 $D=0
M904 6 169 171 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=25000 $D=0
M905 7 170 172 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=29630 $D=0
M906 173 1 4 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=25000 $D=0
M907 174 1 4 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=29630 $D=0
M908 5 169 173 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=25000 $D=0
M909 5 170 174 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=29630 $D=0
M910 175 1 6 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=25000 $D=0
M911 176 1 7 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=29630 $D=0
M912 6 169 175 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=25000 $D=0
M913 7 170 176 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=29630 $D=0
M914 179 9 175 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=25000 $D=0
M915 180 9 176 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=29630 $D=0
M916 177 9 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=25000 $D=0
M917 178 9 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=29630 $D=0
M918 181 9 173 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=25000 $D=0
M919 182 9 174 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=29630 $D=0
M920 171 177 181 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=25000 $D=0
M921 172 178 182 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=29630 $D=0
M922 183 10 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=25000 $D=0
M923 184 10 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=29630 $D=0
M924 185 10 181 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=25000 $D=0
M925 186 10 182 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=29630 $D=0
M926 179 183 185 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=25000 $D=0
M927 180 184 186 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=29630 $D=0
M928 187 11 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=25000 $D=0
M929 188 11 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=29630 $D=0
M930 189 11 6 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=25000 $D=0
M931 190 11 7 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=29630 $D=0
M932 12 187 189 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=25000 $D=0
M933 13 188 190 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=29630 $D=0
M934 191 11 14 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=25000 $D=0
M935 192 11 15 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=29630 $D=0
M936 193 187 191 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=25000 $D=0
M937 194 188 192 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=29630 $D=0
M938 197 11 195 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=25000 $D=0
M939 198 11 196 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=29630 $D=0
M940 185 187 197 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=25000 $D=0
M941 186 188 198 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=29630 $D=0
M942 201 16 197 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=25000 $D=0
M943 202 16 198 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=29630 $D=0
M944 199 16 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=25000 $D=0
M945 200 16 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=29630 $D=0
M946 203 16 191 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=25000 $D=0
M947 204 16 192 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=29630 $D=0
M948 189 199 203 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=25000 $D=0
M949 190 200 204 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=29630 $D=0
M950 205 17 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=25000 $D=0
M951 206 17 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=29630 $D=0
M952 207 17 203 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=25000 $D=0
M953 208 17 204 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=29630 $D=0
M954 201 205 207 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=25000 $D=0
M955 202 206 208 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=29630 $D=0
M956 164 18 209 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=25000 $D=0
M957 165 18 210 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=29630 $D=0
M958 211 19 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=25000 $D=0
M959 212 19 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=29630 $D=0
M960 213 209 207 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=25000 $D=0
M961 214 210 208 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=29630 $D=0
M962 164 213 684 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=25000 $D=0
M963 165 214 685 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=29630 $D=0
M964 215 684 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=25000 $D=0
M965 216 685 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=29630 $D=0
M966 213 18 215 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=25000 $D=0
M967 214 18 216 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=29630 $D=0
M968 215 211 217 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=25000 $D=0
M969 216 212 218 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=29630 $D=0
M970 221 219 215 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=25000 $D=0
M971 222 220 216 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=29630 $D=0
M972 219 20 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=25000 $D=0
M973 220 20 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=29630 $D=0
M974 164 21 223 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=25000 $D=0
M975 165 21 224 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=29630 $D=0
M976 225 22 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=25000 $D=0
M977 226 22 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=29630 $D=0
M978 227 223 207 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=25000 $D=0
M979 228 224 208 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=29630 $D=0
M980 164 227 686 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=25000 $D=0
M981 165 228 687 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=29630 $D=0
M982 229 686 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=25000 $D=0
M983 230 687 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=29630 $D=0
M984 227 21 229 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=25000 $D=0
M985 228 21 230 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=29630 $D=0
M986 229 225 217 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=25000 $D=0
M987 230 226 218 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=29630 $D=0
M988 221 231 229 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=25000 $D=0
M989 222 232 230 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=29630 $D=0
M990 231 23 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=25000 $D=0
M991 232 23 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=29630 $D=0
M992 164 24 233 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=25000 $D=0
M993 165 24 234 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=29630 $D=0
M994 235 25 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=25000 $D=0
M995 236 25 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=29630 $D=0
M996 237 233 207 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=25000 $D=0
M997 238 234 208 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=29630 $D=0
M998 164 237 688 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=25000 $D=0
M999 165 238 689 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=29630 $D=0
M1000 239 688 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=25000 $D=0
M1001 240 689 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=29630 $D=0
M1002 237 24 239 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=25000 $D=0
M1003 238 24 240 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=29630 $D=0
M1004 239 235 217 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=25000 $D=0
M1005 240 236 218 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=29630 $D=0
M1006 221 241 239 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=25000 $D=0
M1007 222 242 240 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=29630 $D=0
M1008 241 26 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=25000 $D=0
M1009 242 26 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=29630 $D=0
M1010 164 27 243 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=25000 $D=0
M1011 165 27 244 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=29630 $D=0
M1012 245 28 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=25000 $D=0
M1013 246 28 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=29630 $D=0
M1014 247 243 207 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=25000 $D=0
M1015 248 244 208 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=29630 $D=0
M1016 164 247 690 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=25000 $D=0
M1017 165 248 691 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=29630 $D=0
M1018 249 690 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=25000 $D=0
M1019 250 691 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=29630 $D=0
M1020 247 27 249 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=25000 $D=0
M1021 248 27 250 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=29630 $D=0
M1022 249 245 217 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=25000 $D=0
M1023 250 246 218 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=29630 $D=0
M1024 221 251 249 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=25000 $D=0
M1025 222 252 250 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=29630 $D=0
M1026 251 29 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=25000 $D=0
M1027 252 29 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=29630 $D=0
M1028 164 30 253 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=25000 $D=0
M1029 165 30 254 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=29630 $D=0
M1030 255 31 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=25000 $D=0
M1031 256 31 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=29630 $D=0
M1032 257 253 207 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=25000 $D=0
M1033 258 254 208 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=29630 $D=0
M1034 164 257 692 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=25000 $D=0
M1035 165 258 693 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=29630 $D=0
M1036 259 692 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=25000 $D=0
M1037 260 693 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=29630 $D=0
M1038 257 30 259 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=25000 $D=0
M1039 258 30 260 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=29630 $D=0
M1040 259 255 217 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=25000 $D=0
M1041 260 256 218 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=29630 $D=0
M1042 221 261 259 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=25000 $D=0
M1043 222 262 260 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=29630 $D=0
M1044 261 32 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=25000 $D=0
M1045 262 32 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=29630 $D=0
M1046 164 33 263 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=25000 $D=0
M1047 165 33 264 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=29630 $D=0
M1048 265 34 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=25000 $D=0
M1049 266 34 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=29630 $D=0
M1050 267 263 207 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=25000 $D=0
M1051 268 264 208 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=29630 $D=0
M1052 164 267 694 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=25000 $D=0
M1053 165 268 695 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=29630 $D=0
M1054 269 694 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=25000 $D=0
M1055 270 695 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=29630 $D=0
M1056 267 33 269 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=25000 $D=0
M1057 268 33 270 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=29630 $D=0
M1058 269 265 217 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=25000 $D=0
M1059 270 266 218 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=29630 $D=0
M1060 221 271 269 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=25000 $D=0
M1061 222 272 270 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=29630 $D=0
M1062 271 35 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=25000 $D=0
M1063 272 35 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=29630 $D=0
M1064 164 36 273 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=25000 $D=0
M1065 165 36 274 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=29630 $D=0
M1066 275 37 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=25000 $D=0
M1067 276 37 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=29630 $D=0
M1068 277 273 207 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=25000 $D=0
M1069 278 274 208 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=29630 $D=0
M1070 164 277 696 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=25000 $D=0
M1071 165 278 697 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=29630 $D=0
M1072 279 696 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=25000 $D=0
M1073 280 697 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=29630 $D=0
M1074 277 36 279 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=25000 $D=0
M1075 278 36 280 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=29630 $D=0
M1076 279 275 217 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=25000 $D=0
M1077 280 276 218 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=29630 $D=0
M1078 221 281 279 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=25000 $D=0
M1079 222 282 280 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=29630 $D=0
M1080 281 38 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=25000 $D=0
M1081 282 38 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=29630 $D=0
M1082 164 39 283 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=25000 $D=0
M1083 165 39 284 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=29630 $D=0
M1084 285 40 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=25000 $D=0
M1085 286 40 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=29630 $D=0
M1086 287 283 207 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=25000 $D=0
M1087 288 284 208 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=29630 $D=0
M1088 164 287 698 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=25000 $D=0
M1089 165 288 699 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=29630 $D=0
M1090 289 698 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=25000 $D=0
M1091 290 699 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=29630 $D=0
M1092 287 39 289 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=25000 $D=0
M1093 288 39 290 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=29630 $D=0
M1094 289 285 217 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=25000 $D=0
M1095 290 286 218 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=29630 $D=0
M1096 221 291 289 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=25000 $D=0
M1097 222 292 290 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=29630 $D=0
M1098 291 41 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=25000 $D=0
M1099 292 41 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=29630 $D=0
M1100 164 42 293 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=25000 $D=0
M1101 165 42 294 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=29630 $D=0
M1102 295 43 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=25000 $D=0
M1103 296 43 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=29630 $D=0
M1104 297 293 207 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=25000 $D=0
M1105 298 294 208 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=29630 $D=0
M1106 164 297 700 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=25000 $D=0
M1107 165 298 701 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=29630 $D=0
M1108 299 700 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=25000 $D=0
M1109 300 701 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=29630 $D=0
M1110 297 42 299 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=25000 $D=0
M1111 298 42 300 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=29630 $D=0
M1112 299 295 217 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=25000 $D=0
M1113 300 296 218 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=29630 $D=0
M1114 221 301 299 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=25000 $D=0
M1115 222 302 300 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=29630 $D=0
M1116 301 44 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=25000 $D=0
M1117 302 44 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=29630 $D=0
M1118 164 45 303 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=25000 $D=0
M1119 165 45 304 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=29630 $D=0
M1120 305 46 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=25000 $D=0
M1121 306 46 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=29630 $D=0
M1122 307 303 207 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=25000 $D=0
M1123 308 304 208 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=29630 $D=0
M1124 164 307 702 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=25000 $D=0
M1125 165 308 703 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=29630 $D=0
M1126 309 702 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=25000 $D=0
M1127 310 703 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=29630 $D=0
M1128 307 45 309 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=25000 $D=0
M1129 308 45 310 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=29630 $D=0
M1130 309 305 217 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=25000 $D=0
M1131 310 306 218 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=29630 $D=0
M1132 221 311 309 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=25000 $D=0
M1133 222 312 310 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=29630 $D=0
M1134 311 47 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=25000 $D=0
M1135 312 47 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=29630 $D=0
M1136 164 48 313 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=25000 $D=0
M1137 165 48 314 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=29630 $D=0
M1138 315 49 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=25000 $D=0
M1139 316 49 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=29630 $D=0
M1140 317 313 207 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=25000 $D=0
M1141 318 314 208 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=29630 $D=0
M1142 164 317 704 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=25000 $D=0
M1143 165 318 705 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=29630 $D=0
M1144 319 704 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=25000 $D=0
M1145 320 705 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=29630 $D=0
M1146 317 48 319 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=25000 $D=0
M1147 318 48 320 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=29630 $D=0
M1148 319 315 217 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=25000 $D=0
M1149 320 316 218 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=29630 $D=0
M1150 221 321 319 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=25000 $D=0
M1151 222 322 320 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=29630 $D=0
M1152 321 50 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=25000 $D=0
M1153 322 50 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=29630 $D=0
M1154 164 51 323 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=25000 $D=0
M1155 165 51 324 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=29630 $D=0
M1156 325 52 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=25000 $D=0
M1157 326 52 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=29630 $D=0
M1158 327 323 207 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=25000 $D=0
M1159 328 324 208 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=29630 $D=0
M1160 164 327 706 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=25000 $D=0
M1161 165 328 707 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=29630 $D=0
M1162 329 706 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=25000 $D=0
M1163 330 707 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=29630 $D=0
M1164 327 51 329 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=25000 $D=0
M1165 328 51 330 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=29630 $D=0
M1166 329 325 217 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=25000 $D=0
M1167 330 326 218 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=29630 $D=0
M1168 221 331 329 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=25000 $D=0
M1169 222 332 330 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=29630 $D=0
M1170 331 53 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=25000 $D=0
M1171 332 53 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=29630 $D=0
M1172 164 54 333 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=25000 $D=0
M1173 165 54 334 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=29630 $D=0
M1174 335 55 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=25000 $D=0
M1175 336 55 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=29630 $D=0
M1176 337 333 207 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=25000 $D=0
M1177 338 334 208 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=29630 $D=0
M1178 164 337 708 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=25000 $D=0
M1179 165 338 709 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=29630 $D=0
M1180 339 708 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=25000 $D=0
M1181 340 709 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=29630 $D=0
M1182 337 54 339 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=25000 $D=0
M1183 338 54 340 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=29630 $D=0
M1184 339 335 217 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=25000 $D=0
M1185 340 336 218 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=29630 $D=0
M1186 221 341 339 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=25000 $D=0
M1187 222 342 340 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=29630 $D=0
M1188 341 56 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=25000 $D=0
M1189 342 56 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=29630 $D=0
M1190 164 57 343 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=25000 $D=0
M1191 165 57 344 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=29630 $D=0
M1192 345 58 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=25000 $D=0
M1193 346 58 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=29630 $D=0
M1194 347 343 207 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=25000 $D=0
M1195 348 344 208 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=29630 $D=0
M1196 164 347 710 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=25000 $D=0
M1197 165 348 711 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=29630 $D=0
M1198 349 710 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=25000 $D=0
M1199 350 711 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=29630 $D=0
M1200 347 57 349 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=25000 $D=0
M1201 348 57 350 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=29630 $D=0
M1202 349 345 217 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=25000 $D=0
M1203 350 346 218 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=29630 $D=0
M1204 221 351 349 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=25000 $D=0
M1205 222 352 350 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=29630 $D=0
M1206 351 59 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=25000 $D=0
M1207 352 59 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=29630 $D=0
M1208 164 60 353 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=25000 $D=0
M1209 165 60 354 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=29630 $D=0
M1210 355 61 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=25000 $D=0
M1211 356 61 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=29630 $D=0
M1212 357 353 207 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=25000 $D=0
M1213 358 354 208 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=29630 $D=0
M1214 164 357 712 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=25000 $D=0
M1215 165 358 713 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=29630 $D=0
M1216 359 712 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=25000 $D=0
M1217 360 713 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=29630 $D=0
M1218 357 60 359 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=25000 $D=0
M1219 358 60 360 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=29630 $D=0
M1220 359 355 217 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=25000 $D=0
M1221 360 356 218 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=29630 $D=0
M1222 221 361 359 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=25000 $D=0
M1223 222 362 360 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=29630 $D=0
M1224 361 62 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=25000 $D=0
M1225 362 62 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=29630 $D=0
M1226 164 63 363 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=25000 $D=0
M1227 165 63 364 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=29630 $D=0
M1228 365 64 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=25000 $D=0
M1229 366 64 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=29630 $D=0
M1230 367 363 207 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=25000 $D=0
M1231 368 364 208 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=29630 $D=0
M1232 164 367 714 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=25000 $D=0
M1233 165 368 715 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=29630 $D=0
M1234 369 714 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=25000 $D=0
M1235 370 715 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=29630 $D=0
M1236 367 63 369 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=25000 $D=0
M1237 368 63 370 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=29630 $D=0
M1238 369 365 217 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=25000 $D=0
M1239 370 366 218 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=29630 $D=0
M1240 221 371 369 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=25000 $D=0
M1241 222 372 370 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=29630 $D=0
M1242 371 65 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=25000 $D=0
M1243 372 65 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=29630 $D=0
M1244 164 66 373 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=25000 $D=0
M1245 165 66 374 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=29630 $D=0
M1246 375 67 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=25000 $D=0
M1247 376 67 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=29630 $D=0
M1248 377 373 207 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=25000 $D=0
M1249 378 374 208 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=29630 $D=0
M1250 164 377 716 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=25000 $D=0
M1251 165 378 717 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=29630 $D=0
M1252 379 716 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=25000 $D=0
M1253 380 717 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=29630 $D=0
M1254 377 66 379 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=25000 $D=0
M1255 378 66 380 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=29630 $D=0
M1256 379 375 217 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=25000 $D=0
M1257 380 376 218 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=29630 $D=0
M1258 221 381 379 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=25000 $D=0
M1259 222 382 380 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=29630 $D=0
M1260 381 68 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=25000 $D=0
M1261 382 68 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=29630 $D=0
M1262 164 69 383 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=25000 $D=0
M1263 165 69 384 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=29630 $D=0
M1264 385 70 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=25000 $D=0
M1265 386 70 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=29630 $D=0
M1266 387 383 207 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=25000 $D=0
M1267 388 384 208 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=29630 $D=0
M1268 164 387 718 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=25000 $D=0
M1269 165 388 719 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=29630 $D=0
M1270 389 718 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=25000 $D=0
M1271 390 719 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=29630 $D=0
M1272 387 69 389 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=25000 $D=0
M1273 388 69 390 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=29630 $D=0
M1274 389 385 217 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=25000 $D=0
M1275 390 386 218 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=29630 $D=0
M1276 221 391 389 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=25000 $D=0
M1277 222 392 390 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=29630 $D=0
M1278 391 71 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=25000 $D=0
M1279 392 71 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=29630 $D=0
M1280 164 72 393 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=25000 $D=0
M1281 165 72 394 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=29630 $D=0
M1282 395 73 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=25000 $D=0
M1283 396 73 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=29630 $D=0
M1284 397 393 207 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=25000 $D=0
M1285 398 394 208 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=29630 $D=0
M1286 164 397 720 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=25000 $D=0
M1287 165 398 721 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=29630 $D=0
M1288 399 720 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=25000 $D=0
M1289 400 721 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=29630 $D=0
M1290 397 72 399 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=25000 $D=0
M1291 398 72 400 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=29630 $D=0
M1292 399 395 217 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=25000 $D=0
M1293 400 396 218 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=29630 $D=0
M1294 221 401 399 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=25000 $D=0
M1295 222 402 400 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=29630 $D=0
M1296 401 74 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=25000 $D=0
M1297 402 74 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=29630 $D=0
M1298 164 75 403 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=25000 $D=0
M1299 165 75 404 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=29630 $D=0
M1300 405 76 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=25000 $D=0
M1301 406 76 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=29630 $D=0
M1302 407 403 207 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=25000 $D=0
M1303 408 404 208 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=29630 $D=0
M1304 164 407 722 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=25000 $D=0
M1305 165 408 723 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=29630 $D=0
M1306 409 722 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=25000 $D=0
M1307 410 723 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=29630 $D=0
M1308 407 75 409 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=25000 $D=0
M1309 408 75 410 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=29630 $D=0
M1310 409 405 217 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=25000 $D=0
M1311 410 406 218 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=29630 $D=0
M1312 221 411 409 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=25000 $D=0
M1313 222 412 410 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=29630 $D=0
M1314 411 77 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=25000 $D=0
M1315 412 77 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=29630 $D=0
M1316 164 78 413 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=25000 $D=0
M1317 165 78 414 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=29630 $D=0
M1318 415 79 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=25000 $D=0
M1319 416 79 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=29630 $D=0
M1320 417 413 207 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=25000 $D=0
M1321 418 414 208 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=29630 $D=0
M1322 164 417 724 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=25000 $D=0
M1323 165 418 725 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=29630 $D=0
M1324 419 724 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=25000 $D=0
M1325 420 725 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=29630 $D=0
M1326 417 78 419 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=25000 $D=0
M1327 418 78 420 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=29630 $D=0
M1328 419 415 217 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=25000 $D=0
M1329 420 416 218 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=29630 $D=0
M1330 221 421 419 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=25000 $D=0
M1331 222 422 420 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=29630 $D=0
M1332 421 80 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=25000 $D=0
M1333 422 80 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=29630 $D=0
M1334 164 81 423 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=25000 $D=0
M1335 165 81 424 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=29630 $D=0
M1336 425 82 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=25000 $D=0
M1337 426 82 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=29630 $D=0
M1338 427 423 207 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=25000 $D=0
M1339 428 424 208 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=29630 $D=0
M1340 164 427 726 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=25000 $D=0
M1341 165 428 727 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=29630 $D=0
M1342 429 726 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=25000 $D=0
M1343 430 727 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=29630 $D=0
M1344 427 81 429 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=25000 $D=0
M1345 428 81 430 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=29630 $D=0
M1346 429 425 217 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=25000 $D=0
M1347 430 426 218 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=29630 $D=0
M1348 221 431 429 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=25000 $D=0
M1349 222 432 430 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=29630 $D=0
M1350 431 83 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=25000 $D=0
M1351 432 83 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=29630 $D=0
M1352 164 84 433 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=25000 $D=0
M1353 165 84 434 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=29630 $D=0
M1354 435 85 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=25000 $D=0
M1355 436 85 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=29630 $D=0
M1356 437 433 207 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=25000 $D=0
M1357 438 434 208 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=29630 $D=0
M1358 164 437 728 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=25000 $D=0
M1359 165 438 729 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=29630 $D=0
M1360 439 728 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=25000 $D=0
M1361 440 729 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=29630 $D=0
M1362 437 84 439 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=25000 $D=0
M1363 438 84 440 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=29630 $D=0
M1364 439 435 217 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=25000 $D=0
M1365 440 436 218 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=29630 $D=0
M1366 221 441 439 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=25000 $D=0
M1367 222 442 440 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=29630 $D=0
M1368 441 86 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=25000 $D=0
M1369 442 86 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=29630 $D=0
M1370 164 87 443 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=25000 $D=0
M1371 165 87 444 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=29630 $D=0
M1372 445 88 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=25000 $D=0
M1373 446 88 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=29630 $D=0
M1374 447 443 207 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=25000 $D=0
M1375 448 444 208 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=29630 $D=0
M1376 164 447 730 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=25000 $D=0
M1377 165 448 731 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=29630 $D=0
M1378 449 730 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=25000 $D=0
M1379 450 731 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=29630 $D=0
M1380 447 87 449 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=25000 $D=0
M1381 448 87 450 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=29630 $D=0
M1382 449 445 217 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=25000 $D=0
M1383 450 446 218 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=29630 $D=0
M1384 221 451 449 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=25000 $D=0
M1385 222 452 450 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=29630 $D=0
M1386 451 89 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=25000 $D=0
M1387 452 89 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=29630 $D=0
M1388 164 90 453 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=25000 $D=0
M1389 165 90 454 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=29630 $D=0
M1390 455 91 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=25000 $D=0
M1391 456 91 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=29630 $D=0
M1392 457 453 207 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=25000 $D=0
M1393 458 454 208 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=29630 $D=0
M1394 164 457 732 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=25000 $D=0
M1395 165 458 733 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=29630 $D=0
M1396 459 732 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=25000 $D=0
M1397 460 733 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=29630 $D=0
M1398 457 90 459 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=25000 $D=0
M1399 458 90 460 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=29630 $D=0
M1400 459 455 217 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=25000 $D=0
M1401 460 456 218 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=29630 $D=0
M1402 221 461 459 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=25000 $D=0
M1403 222 462 460 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=29630 $D=0
M1404 461 92 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=25000 $D=0
M1405 462 92 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=29630 $D=0
M1406 164 93 463 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=25000 $D=0
M1407 165 93 464 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=29630 $D=0
M1408 465 94 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=25000 $D=0
M1409 466 94 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=29630 $D=0
M1410 467 463 207 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=25000 $D=0
M1411 468 464 208 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=29630 $D=0
M1412 164 467 734 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=25000 $D=0
M1413 165 468 735 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=29630 $D=0
M1414 469 734 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=25000 $D=0
M1415 470 735 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=29630 $D=0
M1416 467 93 469 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=25000 $D=0
M1417 468 93 470 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=29630 $D=0
M1418 469 465 217 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=25000 $D=0
M1419 470 466 218 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=29630 $D=0
M1420 221 471 469 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=25000 $D=0
M1421 222 472 470 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=29630 $D=0
M1422 471 95 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=25000 $D=0
M1423 472 95 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=29630 $D=0
M1424 164 96 473 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=25000 $D=0
M1425 165 96 474 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=29630 $D=0
M1426 475 97 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=25000 $D=0
M1427 476 97 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=29630 $D=0
M1428 477 473 207 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=25000 $D=0
M1429 478 474 208 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=29630 $D=0
M1430 164 477 736 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=25000 $D=0
M1431 165 478 737 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=29630 $D=0
M1432 479 736 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=25000 $D=0
M1433 480 737 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=29630 $D=0
M1434 477 96 479 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=25000 $D=0
M1435 478 96 480 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=29630 $D=0
M1436 479 475 217 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=25000 $D=0
M1437 480 476 218 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=29630 $D=0
M1438 221 481 479 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=25000 $D=0
M1439 222 482 480 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=29630 $D=0
M1440 481 98 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=25000 $D=0
M1441 482 98 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=29630 $D=0
M1442 164 99 483 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=25000 $D=0
M1443 165 99 484 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=29630 $D=0
M1444 485 100 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=25000 $D=0
M1445 486 100 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=29630 $D=0
M1446 487 483 207 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=25000 $D=0
M1447 488 484 208 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=29630 $D=0
M1448 164 487 738 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=25000 $D=0
M1449 165 488 739 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=29630 $D=0
M1450 489 738 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=25000 $D=0
M1451 490 739 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=29630 $D=0
M1452 487 99 489 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=25000 $D=0
M1453 488 99 490 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=29630 $D=0
M1454 489 485 217 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=25000 $D=0
M1455 490 486 218 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=29630 $D=0
M1456 221 491 489 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=25000 $D=0
M1457 222 492 490 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=29630 $D=0
M1458 491 101 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=25000 $D=0
M1459 492 101 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=29630 $D=0
M1460 164 102 493 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=25000 $D=0
M1461 165 102 494 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=29630 $D=0
M1462 495 103 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=25000 $D=0
M1463 496 103 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=29630 $D=0
M1464 497 493 207 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=25000 $D=0
M1465 498 494 208 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=29630 $D=0
M1466 164 497 740 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=25000 $D=0
M1467 165 498 741 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=29630 $D=0
M1468 499 740 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=25000 $D=0
M1469 500 741 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=29630 $D=0
M1470 497 102 499 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=25000 $D=0
M1471 498 102 500 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=29630 $D=0
M1472 499 495 217 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=25000 $D=0
M1473 500 496 218 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=29630 $D=0
M1474 221 501 499 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=25000 $D=0
M1475 222 502 500 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=29630 $D=0
M1476 501 104 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=25000 $D=0
M1477 502 104 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=29630 $D=0
M1478 164 105 503 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=25000 $D=0
M1479 165 105 504 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=29630 $D=0
M1480 505 106 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=25000 $D=0
M1481 506 106 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=29630 $D=0
M1482 507 503 207 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=25000 $D=0
M1483 508 504 208 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=29630 $D=0
M1484 164 507 742 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=25000 $D=0
M1485 165 508 743 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=29630 $D=0
M1486 509 742 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=25000 $D=0
M1487 510 743 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=29630 $D=0
M1488 507 105 509 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=25000 $D=0
M1489 508 105 510 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=29630 $D=0
M1490 509 505 217 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=25000 $D=0
M1491 510 506 218 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=29630 $D=0
M1492 221 511 509 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=25000 $D=0
M1493 222 512 510 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=29630 $D=0
M1494 511 107 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=25000 $D=0
M1495 512 107 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=29630 $D=0
M1496 164 108 513 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=25000 $D=0
M1497 165 108 514 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=29630 $D=0
M1498 515 109 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=25000 $D=0
M1499 516 109 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=29630 $D=0
M1500 517 513 207 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=25000 $D=0
M1501 518 514 208 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=29630 $D=0
M1502 164 517 744 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=25000 $D=0
M1503 165 518 745 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=29630 $D=0
M1504 519 744 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=25000 $D=0
M1505 520 745 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=29630 $D=0
M1506 517 108 519 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=25000 $D=0
M1507 518 108 520 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=29630 $D=0
M1508 519 515 217 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=25000 $D=0
M1509 520 516 218 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=29630 $D=0
M1510 221 521 519 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=25000 $D=0
M1511 222 522 520 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=29630 $D=0
M1512 521 110 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=25000 $D=0
M1513 522 110 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=29630 $D=0
M1514 164 111 523 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=25000 $D=0
M1515 165 111 524 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=29630 $D=0
M1516 525 112 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=25000 $D=0
M1517 526 112 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=29630 $D=0
M1518 6 525 217 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=25000 $D=0
M1519 7 526 218 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=29630 $D=0
M1520 221 523 6 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=25000 $D=0
M1521 222 524 7 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=29630 $D=0
M1522 164 529 527 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=25000 $D=0
M1523 165 530 528 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=29630 $D=0
M1524 529 113 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=25000 $D=0
M1525 530 113 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=29630 $D=0
M1526 746 217 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=25000 $D=0
M1527 747 218 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=29630 $D=0
M1528 531 529 746 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=25000 $D=0
M1529 532 530 747 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=29630 $D=0
M1530 164 531 533 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=25000 $D=0
M1531 165 532 534 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=29630 $D=0
M1532 748 533 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=25000 $D=0
M1533 749 534 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=29630 $D=0
M1534 531 527 748 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=25000 $D=0
M1535 532 528 749 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=29630 $D=0
M1536 164 537 535 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=25000 $D=0
M1537 165 538 536 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=29630 $D=0
M1538 537 113 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=25000 $D=0
M1539 538 113 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=29630 $D=0
M1540 750 221 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=25000 $D=0
M1541 751 222 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=29630 $D=0
M1542 539 537 750 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=25000 $D=0
M1543 540 538 751 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=29630 $D=0
M1544 164 539 114 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=25000 $D=0
M1545 165 540 115 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=29630 $D=0
M1546 752 114 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=25000 $D=0
M1547 753 115 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=29630 $D=0
M1548 539 535 752 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=25000 $D=0
M1549 540 536 753 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=29630 $D=0
M1550 541 116 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=25000 $D=0
M1551 542 116 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=29630 $D=0
M1552 543 116 533 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=25000 $D=0
M1553 544 116 534 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=29630 $D=0
M1554 117 541 543 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=25000 $D=0
M1555 118 542 544 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=29630 $D=0
M1556 545 119 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=25000 $D=0
M1557 546 119 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=29630 $D=0
M1558 547 119 114 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=25000 $D=0
M1559 548 119 115 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=29630 $D=0
M1560 754 545 547 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=25000 $D=0
M1561 755 546 548 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=29630 $D=0
M1562 164 114 754 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=25000 $D=0
M1563 165 115 755 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=29630 $D=0
M1564 549 120 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=25000 $D=0
M1565 550 120 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=29630 $D=0
M1566 551 120 547 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=25000 $D=0
M1567 552 120 548 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=29630 $D=0
M1568 12 549 551 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=25000 $D=0
M1569 13 550 552 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=29630 $D=0
M1570 555 553 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=25000 $D=0
M1571 556 554 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=29630 $D=0
M1572 164 559 557 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=25000 $D=0
M1573 165 560 558 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=29630 $D=0
M1574 561 543 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=25000 $D=0
M1575 562 544 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=29630 $D=0
M1576 559 543 553 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=25000 $D=0
M1577 560 544 554 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=29630 $D=0
M1578 555 561 559 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=25000 $D=0
M1579 556 562 560 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=29630 $D=0
M1580 563 557 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=25000 $D=0
M1581 564 558 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=29630 $D=0
M1582 121 557 551 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=25000 $D=0
M1583 553 558 552 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=29630 $D=0
M1584 543 563 121 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=25000 $D=0
M1585 544 564 553 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=29630 $D=0
M1586 565 121 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=25000 $D=0
M1587 566 553 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=29630 $D=0
M1588 567 557 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=25000 $D=0
M1589 568 558 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=29630 $D=0
M1590 569 557 565 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=25000 $D=0
M1591 570 558 566 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=29630 $D=0
M1592 551 567 569 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=25000 $D=0
M1593 552 568 570 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=29630 $D=0
M1594 774 543 164 164 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=24640 $D=0
M1595 775 544 165 165 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=29270 $D=0
M1596 571 551 774 164 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=24640 $D=0
M1597 572 552 775 165 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=29270 $D=0
M1598 573 569 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=25000 $D=0
M1599 574 570 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=29630 $D=0
M1600 575 543 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=25000 $D=0
M1601 576 544 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=29630 $D=0
M1602 164 551 575 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=25000 $D=0
M1603 165 552 576 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=29630 $D=0
M1604 577 543 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=25000 $D=0
M1605 578 544 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=29630 $D=0
M1606 164 551 577 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=25000 $D=0
M1607 165 552 578 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=29630 $D=0
M1608 776 543 164 164 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=24820 $D=0
M1609 777 544 165 165 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=29450 $D=0
M1610 581 551 776 164 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=24820 $D=0
M1611 582 552 777 165 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=29450 $D=0
M1612 164 577 581 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=25000 $D=0
M1613 165 578 582 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=29630 $D=0
M1614 583 126 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=25000 $D=0
M1615 584 126 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=29630 $D=0
M1616 585 126 571 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=25000 $D=0
M1617 586 126 572 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=29630 $D=0
M1618 575 583 585 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=25000 $D=0
M1619 576 584 586 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=29630 $D=0
M1620 587 126 573 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=25000 $D=0
M1621 588 126 574 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=29630 $D=0
M1622 581 583 587 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=25000 $D=0
M1623 582 584 588 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=29630 $D=0
M1624 589 127 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=25000 $D=0
M1625 590 127 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=29630 $D=0
M1626 591 127 587 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=25000 $D=0
M1627 592 127 588 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=29630 $D=0
M1628 585 589 591 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=25000 $D=0
M1629 586 590 592 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=29630 $D=0
M1630 14 591 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=25000 $D=0
M1631 15 592 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=29630 $D=0
M1632 593 128 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=25000 $D=0
M1633 594 128 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=29630 $D=0
M1634 595 128 129 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=25000 $D=0
M1635 596 128 130 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=29630 $D=0
M1636 131 593 595 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=25000 $D=0
M1637 132 594 596 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=29630 $D=0
M1638 597 128 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=25000 $D=0
M1639 598 128 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=29630 $D=0
M1640 600 128 133 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=25000 $D=0
M1641 601 128 135 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=29630 $D=0
M1642 136 597 600 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=25000 $D=0
M1643 134 598 601 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=29630 $D=0
M1644 602 128 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=25000 $D=0
M1645 603 128 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=29630 $D=0
M1646 604 128 125 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=25000 $D=0
M1647 605 128 124 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=29630 $D=0
M1648 137 602 604 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=25000 $D=0
M1649 138 603 605 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=29630 $D=0
M1650 606 128 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=25000 $D=0
M1651 607 128 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=29630 $D=0
M1652 608 128 139 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=25000 $D=0
M1653 609 128 140 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=29630 $D=0
M1654 141 606 608 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=25000 $D=0
M1655 141 607 609 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=29630 $D=0
M1656 610 128 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=25000 $D=0
M1657 611 128 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=29630 $D=0
M1658 612 128 142 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=25000 $D=0
M1659 613 128 143 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=29630 $D=0
M1660 141 610 612 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=25000 $D=0
M1661 141 611 613 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=29630 $D=0
M1662 164 543 764 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=25000 $D=0
M1663 165 544 765 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=29630 $D=0
M1664 132 764 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=25000 $D=0
M1665 129 765 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=29630 $D=0
M1666 614 144 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=25000 $D=0
M1667 615 144 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=29630 $D=0
M1668 145 144 132 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=25000 $D=0
M1669 146 144 129 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=29630 $D=0
M1670 595 614 145 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=25000 $D=0
M1671 596 615 146 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=29630 $D=0
M1672 616 147 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=25000 $D=0
M1673 617 147 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=29630 $D=0
M1674 148 147 145 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=25000 $D=0
M1675 123 147 146 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=29630 $D=0
M1676 600 616 148 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=25000 $D=0
M1677 601 617 123 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=29630 $D=0
M1678 618 149 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=25000 $D=0
M1679 619 149 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=29630 $D=0
M1680 150 149 148 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=25000 $D=0
M1681 151 149 123 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=29630 $D=0
M1682 604 618 150 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=25000 $D=0
M1683 605 619 151 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=29630 $D=0
M1684 620 152 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=25000 $D=0
M1685 621 152 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=29630 $D=0
M1686 153 152 150 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=25000 $D=0
M1687 154 152 151 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=29630 $D=0
M1688 608 620 153 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=25000 $D=0
M1689 609 621 154 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=29630 $D=0
M1690 622 155 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=25000 $D=0
M1691 623 155 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=29630 $D=0
M1692 193 155 153 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=25000 $D=0
M1693 194 155 154 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=29630 $D=0
M1694 612 622 193 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=25000 $D=0
M1695 613 623 194 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=29630 $D=0
M1696 624 156 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=25000 $D=0
M1697 625 156 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=29630 $D=0
M1698 626 156 114 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=25000 $D=0
M1699 627 156 115 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=29630 $D=0
M1700 12 624 626 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=25000 $D=0
M1701 13 625 627 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=29630 $D=0
M1702 628 533 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=25000 $D=0
M1703 629 534 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=29630 $D=0
M1704 164 626 628 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=25000 $D=0
M1705 165 627 629 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=29630 $D=0
M1706 778 533 164 164 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=24820 $D=0
M1707 779 534 165 165 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=29450 $D=0
M1708 632 626 778 164 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=24820 $D=0
M1709 633 627 779 165 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=29450 $D=0
M1710 164 628 632 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=25000 $D=0
M1711 165 629 633 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=29630 $D=0
M1712 766 157 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=25000 $D=0
M1713 767 634 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=29630 $D=0
M1714 164 632 766 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=25000 $D=0
M1715 165 633 767 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=29630 $D=0
M1716 634 766 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=25000 $D=0
M1717 635 767 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=29630 $D=0
M1718 780 533 164 164 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=24640 $D=0
M1719 781 534 165 165 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=29270 $D=0
M1720 636 638 780 164 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=24640 $D=0
M1721 637 639 781 165 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=29270 $D=0
M1722 638 626 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=25000 $D=0
M1723 639 627 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=29630 $D=0
M1724 640 636 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=25000 $D=0
M1725 641 637 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=29630 $D=0
M1726 164 157 640 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=25000 $D=0
M1727 165 634 641 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=29630 $D=0
M1728 643 158 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=25000 $D=0
M1729 644 642 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=29630 $D=0
M1730 642 640 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=25000 $D=0
M1731 159 641 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=29630 $D=0
M1732 164 643 642 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=25000 $D=0
M1733 165 644 159 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=29630 $D=0
M1734 646 645 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=25000 $D=0
M1735 647 160 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=29630 $D=0
M1736 164 650 648 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=25000 $D=0
M1737 165 651 649 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=29630 $D=0
M1738 652 117 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=25000 $D=0
M1739 653 118 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=29630 $D=0
M1740 650 117 645 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=25000 $D=0
M1741 651 118 160 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=29630 $D=0
M1742 646 652 650 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=25000 $D=0
M1743 647 653 651 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=29630 $D=0
M1744 654 648 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=25000 $D=0
M1745 655 649 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=29630 $D=0
M1746 161 648 6 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=25000 $D=0
M1747 645 649 7 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=29630 $D=0
M1748 117 654 161 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=25000 $D=0
M1749 118 655 645 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=29630 $D=0
M1750 656 161 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=25000 $D=0
M1751 657 645 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=29630 $D=0
M1752 658 648 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=25000 $D=0
M1753 659 649 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=29630 $D=0
M1754 195 648 656 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=25000 $D=0
M1755 196 649 657 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=29630 $D=0
M1756 6 658 195 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=25000 $D=0
M1757 7 659 196 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=29630 $D=0
M1758 660 162 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=25000 $D=0
M1759 661 162 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=29630 $D=0
M1760 662 162 195 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=25000 $D=0
M1761 663 162 196 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=29630 $D=0
M1762 14 660 662 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=25000 $D=0
M1763 15 661 663 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=29630 $D=0
M1764 664 163 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=25000 $D=0
M1765 665 163 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=29630 $D=0
M1766 163 163 662 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=25000 $D=0
M1767 163 163 663 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=29630 $D=0
M1768 6 664 163 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=25000 $D=0
M1769 7 665 163 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=29630 $D=0
M1770 666 113 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=25000 $D=0
M1771 667 113 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=29630 $D=0
M1772 164 666 668 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=25000 $D=0
M1773 165 667 669 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=29630 $D=0
M1774 670 113 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=25000 $D=0
M1775 671 113 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=29630 $D=0
M1776 672 668 163 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=25000 $D=0
M1777 673 669 163 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=29630 $D=0
M1778 164 672 768 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=25000 $D=0
M1779 165 673 769 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=29630 $D=0
M1780 674 768 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=25000 $D=0
M1781 675 769 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=29630 $D=0
M1782 672 666 674 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=25000 $D=0
M1783 673 667 675 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=29630 $D=0
M1784 676 670 674 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=25000 $D=0
M1785 677 671 675 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=29630 $D=0
M1786 164 680 678 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=25000 $D=0
M1787 165 681 679 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=29630 $D=0
M1788 680 113 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=25000 $D=0
M1789 681 113 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=29630 $D=0
M1790 770 676 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=25000 $D=0
M1791 771 677 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=29630 $D=0
M1792 682 680 770 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=25000 $D=0
M1793 683 681 771 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=29630 $D=0
M1794 164 682 117 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=25000 $D=0
M1795 165 683 118 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=29630 $D=0
M1796 772 117 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=25000 $D=0
M1797 773 118 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=29630 $D=0
M1798 682 678 772 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=25000 $D=0
M1799 683 679 773 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=29630 $D=0
.ENDS
***************************************
.SUBCKT ICV_40 1 2 3 4 5 6 7 9 10 11 12 13 14 15 16 17 18 19 20 21
+ 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41
+ 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61
+ 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81
+ 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101
+ 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121
+ 122 123 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141 142
+ 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162
+ 163 164 165
** N=793 EP=163 IP=1514 FDC=1800
M0 169 1 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=14490 $D=1
M1 170 1 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=19120 $D=1
M2 171 169 2 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=14490 $D=1
M3 172 170 3 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=19120 $D=1
M4 6 1 171 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=14490 $D=1
M5 7 1 172 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=19120 $D=1
M6 173 169 4 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=14490 $D=1
M7 174 170 4 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=19120 $D=1
M8 5 1 173 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=14490 $D=1
M9 5 1 174 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=19120 $D=1
M10 175 169 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=14490 $D=1
M11 176 170 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=19120 $D=1
M12 6 1 175 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=14490 $D=1
M13 7 1 176 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=19120 $D=1
M14 179 177 175 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=14490 $D=1
M15 180 178 176 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=19120 $D=1
M16 177 9 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=14490 $D=1
M17 178 9 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=19120 $D=1
M18 181 177 173 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=14490 $D=1
M19 182 178 174 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=19120 $D=1
M20 171 9 181 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=14490 $D=1
M21 172 9 182 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=19120 $D=1
M22 183 10 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=14490 $D=1
M23 184 10 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=19120 $D=1
M24 185 183 181 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=14490 $D=1
M25 186 184 182 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=19120 $D=1
M26 179 10 185 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=14490 $D=1
M27 180 10 186 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=19120 $D=1
M28 187 11 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=14490 $D=1
M29 188 11 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=19120 $D=1
M30 189 187 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=14490 $D=1
M31 190 188 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=19120 $D=1
M32 12 11 189 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=14490 $D=1
M33 13 11 190 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=19120 $D=1
M34 191 187 14 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=14490 $D=1
M35 192 188 15 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=19120 $D=1
M36 193 11 191 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=14490 $D=1
M37 194 11 192 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=19120 $D=1
M38 197 187 195 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=14490 $D=1
M39 198 188 196 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=19120 $D=1
M40 185 11 197 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=14490 $D=1
M41 186 11 198 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=19120 $D=1
M42 201 199 197 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=14490 $D=1
M43 202 200 198 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=19120 $D=1
M44 199 16 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=14490 $D=1
M45 200 16 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=19120 $D=1
M46 203 199 191 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=14490 $D=1
M47 204 200 192 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=19120 $D=1
M48 189 16 203 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=14490 $D=1
M49 190 16 204 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=19120 $D=1
M50 205 17 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=14490 $D=1
M51 206 17 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=19120 $D=1
M52 207 205 203 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=14490 $D=1
M53 208 206 204 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=19120 $D=1
M54 201 17 207 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=14490 $D=1
M55 202 17 208 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=19120 $D=1
M56 6 18 209 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=14490 $D=1
M57 7 18 210 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=19120 $D=1
M58 211 19 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=14490 $D=1
M59 212 19 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=19120 $D=1
M60 213 18 207 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=14490 $D=1
M61 214 18 208 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=19120 $D=1
M62 6 213 684 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=14490 $D=1
M63 7 214 685 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=19120 $D=1
M64 215 684 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=14490 $D=1
M65 216 685 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=19120 $D=1
M66 213 209 215 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=14490 $D=1
M67 214 210 216 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=19120 $D=1
M68 215 19 217 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=14490 $D=1
M69 216 19 218 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=19120 $D=1
M70 221 20 215 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=14490 $D=1
M71 222 20 216 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=19120 $D=1
M72 219 20 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=14490 $D=1
M73 220 20 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=19120 $D=1
M74 6 21 223 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=14490 $D=1
M75 7 21 224 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=19120 $D=1
M76 225 22 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=14490 $D=1
M77 226 22 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=19120 $D=1
M78 227 21 207 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=14490 $D=1
M79 228 21 208 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=19120 $D=1
M80 6 227 686 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=14490 $D=1
M81 7 228 687 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=19120 $D=1
M82 229 686 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=14490 $D=1
M83 230 687 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=19120 $D=1
M84 227 223 229 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=14490 $D=1
M85 228 224 230 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=19120 $D=1
M86 229 22 217 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=14490 $D=1
M87 230 22 218 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=19120 $D=1
M88 221 23 229 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=14490 $D=1
M89 222 23 230 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=19120 $D=1
M90 231 23 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=14490 $D=1
M91 232 23 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=19120 $D=1
M92 6 24 233 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=14490 $D=1
M93 7 24 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=19120 $D=1
M94 235 25 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=14490 $D=1
M95 236 25 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=19120 $D=1
M96 237 24 207 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=14490 $D=1
M97 238 24 208 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=19120 $D=1
M98 6 237 688 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=14490 $D=1
M99 7 238 689 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=19120 $D=1
M100 239 688 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=14490 $D=1
M101 240 689 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=19120 $D=1
M102 237 233 239 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=14490 $D=1
M103 238 234 240 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=19120 $D=1
M104 239 25 217 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=14490 $D=1
M105 240 25 218 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=19120 $D=1
M106 221 26 239 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=14490 $D=1
M107 222 26 240 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=19120 $D=1
M108 241 26 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=14490 $D=1
M109 242 26 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=19120 $D=1
M110 6 27 243 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=14490 $D=1
M111 7 27 244 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=19120 $D=1
M112 245 28 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=14490 $D=1
M113 246 28 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=19120 $D=1
M114 247 27 207 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=14490 $D=1
M115 248 27 208 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=19120 $D=1
M116 6 247 690 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=14490 $D=1
M117 7 248 691 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=19120 $D=1
M118 249 690 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=14490 $D=1
M119 250 691 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=19120 $D=1
M120 247 243 249 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=14490 $D=1
M121 248 244 250 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=19120 $D=1
M122 249 28 217 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=14490 $D=1
M123 250 28 218 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=19120 $D=1
M124 221 29 249 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=14490 $D=1
M125 222 29 250 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=19120 $D=1
M126 251 29 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=14490 $D=1
M127 252 29 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=19120 $D=1
M128 6 30 253 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=14490 $D=1
M129 7 30 254 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=19120 $D=1
M130 255 31 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=14490 $D=1
M131 256 31 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=19120 $D=1
M132 257 30 207 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=14490 $D=1
M133 258 30 208 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=19120 $D=1
M134 6 257 692 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=14490 $D=1
M135 7 258 693 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=19120 $D=1
M136 259 692 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=14490 $D=1
M137 260 693 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=19120 $D=1
M138 257 253 259 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=14490 $D=1
M139 258 254 260 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=19120 $D=1
M140 259 31 217 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=14490 $D=1
M141 260 31 218 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=19120 $D=1
M142 221 32 259 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=14490 $D=1
M143 222 32 260 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=19120 $D=1
M144 261 32 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=14490 $D=1
M145 262 32 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=19120 $D=1
M146 6 33 263 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=14490 $D=1
M147 7 33 264 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=19120 $D=1
M148 265 34 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=14490 $D=1
M149 266 34 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=19120 $D=1
M150 267 33 207 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=14490 $D=1
M151 268 33 208 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=19120 $D=1
M152 6 267 694 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=14490 $D=1
M153 7 268 695 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=19120 $D=1
M154 269 694 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=14490 $D=1
M155 270 695 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=19120 $D=1
M156 267 263 269 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=14490 $D=1
M157 268 264 270 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=19120 $D=1
M158 269 34 217 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=14490 $D=1
M159 270 34 218 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=19120 $D=1
M160 221 35 269 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=14490 $D=1
M161 222 35 270 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=19120 $D=1
M162 271 35 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=14490 $D=1
M163 272 35 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=19120 $D=1
M164 6 36 273 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=14490 $D=1
M165 7 36 274 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=19120 $D=1
M166 275 37 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=14490 $D=1
M167 276 37 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=19120 $D=1
M168 277 36 207 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=14490 $D=1
M169 278 36 208 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=19120 $D=1
M170 6 277 696 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=14490 $D=1
M171 7 278 697 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=19120 $D=1
M172 279 696 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=14490 $D=1
M173 280 697 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=19120 $D=1
M174 277 273 279 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=14490 $D=1
M175 278 274 280 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=19120 $D=1
M176 279 37 217 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=14490 $D=1
M177 280 37 218 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=19120 $D=1
M178 221 38 279 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=14490 $D=1
M179 222 38 280 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=19120 $D=1
M180 281 38 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=14490 $D=1
M181 282 38 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=19120 $D=1
M182 6 39 283 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=14490 $D=1
M183 7 39 284 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=19120 $D=1
M184 285 40 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=14490 $D=1
M185 286 40 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=19120 $D=1
M186 287 39 207 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=14490 $D=1
M187 288 39 208 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=19120 $D=1
M188 6 287 698 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=14490 $D=1
M189 7 288 699 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=19120 $D=1
M190 289 698 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=14490 $D=1
M191 290 699 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=19120 $D=1
M192 287 283 289 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=14490 $D=1
M193 288 284 290 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=19120 $D=1
M194 289 40 217 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=14490 $D=1
M195 290 40 218 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=19120 $D=1
M196 221 41 289 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=14490 $D=1
M197 222 41 290 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=19120 $D=1
M198 291 41 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=14490 $D=1
M199 292 41 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=19120 $D=1
M200 6 42 293 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=14490 $D=1
M201 7 42 294 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=19120 $D=1
M202 295 43 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=14490 $D=1
M203 296 43 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=19120 $D=1
M204 297 42 207 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=14490 $D=1
M205 298 42 208 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=19120 $D=1
M206 6 297 700 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=14490 $D=1
M207 7 298 701 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=19120 $D=1
M208 299 700 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=14490 $D=1
M209 300 701 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=19120 $D=1
M210 297 293 299 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=14490 $D=1
M211 298 294 300 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=19120 $D=1
M212 299 43 217 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=14490 $D=1
M213 300 43 218 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=19120 $D=1
M214 221 44 299 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=14490 $D=1
M215 222 44 300 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=19120 $D=1
M216 301 44 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=14490 $D=1
M217 302 44 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=19120 $D=1
M218 6 45 303 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=14490 $D=1
M219 7 45 304 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=19120 $D=1
M220 305 46 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=14490 $D=1
M221 306 46 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=19120 $D=1
M222 307 45 207 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=14490 $D=1
M223 308 45 208 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=19120 $D=1
M224 6 307 702 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=14490 $D=1
M225 7 308 703 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=19120 $D=1
M226 309 702 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=14490 $D=1
M227 310 703 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=19120 $D=1
M228 307 303 309 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=14490 $D=1
M229 308 304 310 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=19120 $D=1
M230 309 46 217 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=14490 $D=1
M231 310 46 218 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=19120 $D=1
M232 221 47 309 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=14490 $D=1
M233 222 47 310 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=19120 $D=1
M234 311 47 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=14490 $D=1
M235 312 47 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=19120 $D=1
M236 6 48 313 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=14490 $D=1
M237 7 48 314 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=19120 $D=1
M238 315 49 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=14490 $D=1
M239 316 49 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=19120 $D=1
M240 317 48 207 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=14490 $D=1
M241 318 48 208 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=19120 $D=1
M242 6 317 704 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=14490 $D=1
M243 7 318 705 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=19120 $D=1
M244 319 704 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=14490 $D=1
M245 320 705 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=19120 $D=1
M246 317 313 319 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=14490 $D=1
M247 318 314 320 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=19120 $D=1
M248 319 49 217 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=14490 $D=1
M249 320 49 218 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=19120 $D=1
M250 221 50 319 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=14490 $D=1
M251 222 50 320 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=19120 $D=1
M252 321 50 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=14490 $D=1
M253 322 50 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=19120 $D=1
M254 6 51 323 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=14490 $D=1
M255 7 51 324 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=19120 $D=1
M256 325 52 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=14490 $D=1
M257 326 52 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=19120 $D=1
M258 327 51 207 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=14490 $D=1
M259 328 51 208 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=19120 $D=1
M260 6 327 706 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=14490 $D=1
M261 7 328 707 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=19120 $D=1
M262 329 706 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=14490 $D=1
M263 330 707 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=19120 $D=1
M264 327 323 329 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=14490 $D=1
M265 328 324 330 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=19120 $D=1
M266 329 52 217 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=14490 $D=1
M267 330 52 218 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=19120 $D=1
M268 221 53 329 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=14490 $D=1
M269 222 53 330 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=19120 $D=1
M270 331 53 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=14490 $D=1
M271 332 53 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=19120 $D=1
M272 6 54 333 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=14490 $D=1
M273 7 54 334 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=19120 $D=1
M274 335 55 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=14490 $D=1
M275 336 55 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=19120 $D=1
M276 337 54 207 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=14490 $D=1
M277 338 54 208 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=19120 $D=1
M278 6 337 708 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=14490 $D=1
M279 7 338 709 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=19120 $D=1
M280 339 708 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=14490 $D=1
M281 340 709 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=19120 $D=1
M282 337 333 339 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=14490 $D=1
M283 338 334 340 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=19120 $D=1
M284 339 55 217 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=14490 $D=1
M285 340 55 218 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=19120 $D=1
M286 221 56 339 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=14490 $D=1
M287 222 56 340 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=19120 $D=1
M288 341 56 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=14490 $D=1
M289 342 56 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=19120 $D=1
M290 6 57 343 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=14490 $D=1
M291 7 57 344 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=19120 $D=1
M292 345 58 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=14490 $D=1
M293 346 58 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=19120 $D=1
M294 347 57 207 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=14490 $D=1
M295 348 57 208 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=19120 $D=1
M296 6 347 710 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=14490 $D=1
M297 7 348 711 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=19120 $D=1
M298 349 710 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=14490 $D=1
M299 350 711 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=19120 $D=1
M300 347 343 349 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=14490 $D=1
M301 348 344 350 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=19120 $D=1
M302 349 58 217 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=14490 $D=1
M303 350 58 218 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=19120 $D=1
M304 221 59 349 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=14490 $D=1
M305 222 59 350 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=19120 $D=1
M306 351 59 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=14490 $D=1
M307 352 59 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=19120 $D=1
M308 6 60 353 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=14490 $D=1
M309 7 60 354 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=19120 $D=1
M310 355 61 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=14490 $D=1
M311 356 61 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=19120 $D=1
M312 357 60 207 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=14490 $D=1
M313 358 60 208 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=19120 $D=1
M314 6 357 712 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=14490 $D=1
M315 7 358 713 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=19120 $D=1
M316 359 712 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=14490 $D=1
M317 360 713 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=19120 $D=1
M318 357 353 359 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=14490 $D=1
M319 358 354 360 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=19120 $D=1
M320 359 61 217 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=14490 $D=1
M321 360 61 218 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=19120 $D=1
M322 221 62 359 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=14490 $D=1
M323 222 62 360 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=19120 $D=1
M324 361 62 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=14490 $D=1
M325 362 62 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=19120 $D=1
M326 6 63 363 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=14490 $D=1
M327 7 63 364 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=19120 $D=1
M328 365 64 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=14490 $D=1
M329 366 64 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=19120 $D=1
M330 367 63 207 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=14490 $D=1
M331 368 63 208 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=19120 $D=1
M332 6 367 714 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=14490 $D=1
M333 7 368 715 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=19120 $D=1
M334 369 714 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=14490 $D=1
M335 370 715 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=19120 $D=1
M336 367 363 369 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=14490 $D=1
M337 368 364 370 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=19120 $D=1
M338 369 64 217 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=14490 $D=1
M339 370 64 218 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=19120 $D=1
M340 221 65 369 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=14490 $D=1
M341 222 65 370 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=19120 $D=1
M342 371 65 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=14490 $D=1
M343 372 65 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=19120 $D=1
M344 6 66 373 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=14490 $D=1
M345 7 66 374 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=19120 $D=1
M346 375 67 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=14490 $D=1
M347 376 67 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=19120 $D=1
M348 377 66 207 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=14490 $D=1
M349 378 66 208 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=19120 $D=1
M350 6 377 716 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=14490 $D=1
M351 7 378 717 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=19120 $D=1
M352 379 716 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=14490 $D=1
M353 380 717 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=19120 $D=1
M354 377 373 379 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=14490 $D=1
M355 378 374 380 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=19120 $D=1
M356 379 67 217 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=14490 $D=1
M357 380 67 218 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=19120 $D=1
M358 221 68 379 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=14490 $D=1
M359 222 68 380 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=19120 $D=1
M360 381 68 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=14490 $D=1
M361 382 68 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=19120 $D=1
M362 6 69 383 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=14490 $D=1
M363 7 69 384 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=19120 $D=1
M364 385 70 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=14490 $D=1
M365 386 70 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=19120 $D=1
M366 387 69 207 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=14490 $D=1
M367 388 69 208 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=19120 $D=1
M368 6 387 718 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=14490 $D=1
M369 7 388 719 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=19120 $D=1
M370 389 718 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=14490 $D=1
M371 390 719 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=19120 $D=1
M372 387 383 389 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=14490 $D=1
M373 388 384 390 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=19120 $D=1
M374 389 70 217 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=14490 $D=1
M375 390 70 218 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=19120 $D=1
M376 221 71 389 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=14490 $D=1
M377 222 71 390 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=19120 $D=1
M378 391 71 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=14490 $D=1
M379 392 71 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=19120 $D=1
M380 6 72 393 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=14490 $D=1
M381 7 72 394 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=19120 $D=1
M382 395 73 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=14490 $D=1
M383 396 73 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=19120 $D=1
M384 397 72 207 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=14490 $D=1
M385 398 72 208 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=19120 $D=1
M386 6 397 720 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=14490 $D=1
M387 7 398 721 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=19120 $D=1
M388 399 720 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=14490 $D=1
M389 400 721 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=19120 $D=1
M390 397 393 399 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=14490 $D=1
M391 398 394 400 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=19120 $D=1
M392 399 73 217 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=14490 $D=1
M393 400 73 218 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=19120 $D=1
M394 221 74 399 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=14490 $D=1
M395 222 74 400 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=19120 $D=1
M396 401 74 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=14490 $D=1
M397 402 74 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=19120 $D=1
M398 6 75 403 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=14490 $D=1
M399 7 75 404 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=19120 $D=1
M400 405 76 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=14490 $D=1
M401 406 76 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=19120 $D=1
M402 407 75 207 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=14490 $D=1
M403 408 75 208 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=19120 $D=1
M404 6 407 722 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=14490 $D=1
M405 7 408 723 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=19120 $D=1
M406 409 722 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=14490 $D=1
M407 410 723 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=19120 $D=1
M408 407 403 409 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=14490 $D=1
M409 408 404 410 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=19120 $D=1
M410 409 76 217 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=14490 $D=1
M411 410 76 218 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=19120 $D=1
M412 221 77 409 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=14490 $D=1
M413 222 77 410 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=19120 $D=1
M414 411 77 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=14490 $D=1
M415 412 77 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=19120 $D=1
M416 6 78 413 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=14490 $D=1
M417 7 78 414 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=19120 $D=1
M418 415 79 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=14490 $D=1
M419 416 79 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=19120 $D=1
M420 417 78 207 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=14490 $D=1
M421 418 78 208 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=19120 $D=1
M422 6 417 724 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=14490 $D=1
M423 7 418 725 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=19120 $D=1
M424 419 724 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=14490 $D=1
M425 420 725 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=19120 $D=1
M426 417 413 419 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=14490 $D=1
M427 418 414 420 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=19120 $D=1
M428 419 79 217 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=14490 $D=1
M429 420 79 218 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=19120 $D=1
M430 221 80 419 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=14490 $D=1
M431 222 80 420 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=19120 $D=1
M432 421 80 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=14490 $D=1
M433 422 80 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=19120 $D=1
M434 6 81 423 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=14490 $D=1
M435 7 81 424 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=19120 $D=1
M436 425 82 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=14490 $D=1
M437 426 82 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=19120 $D=1
M438 427 81 207 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=14490 $D=1
M439 428 81 208 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=19120 $D=1
M440 6 427 726 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=14490 $D=1
M441 7 428 727 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=19120 $D=1
M442 429 726 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=14490 $D=1
M443 430 727 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=19120 $D=1
M444 427 423 429 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=14490 $D=1
M445 428 424 430 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=19120 $D=1
M446 429 82 217 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=14490 $D=1
M447 430 82 218 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=19120 $D=1
M448 221 83 429 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=14490 $D=1
M449 222 83 430 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=19120 $D=1
M450 431 83 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=14490 $D=1
M451 432 83 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=19120 $D=1
M452 6 84 433 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=14490 $D=1
M453 7 84 434 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=19120 $D=1
M454 435 85 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=14490 $D=1
M455 436 85 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=19120 $D=1
M456 437 84 207 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=14490 $D=1
M457 438 84 208 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=19120 $D=1
M458 6 437 728 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=14490 $D=1
M459 7 438 729 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=19120 $D=1
M460 439 728 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=14490 $D=1
M461 440 729 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=19120 $D=1
M462 437 433 439 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=14490 $D=1
M463 438 434 440 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=19120 $D=1
M464 439 85 217 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=14490 $D=1
M465 440 85 218 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=19120 $D=1
M466 221 86 439 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=14490 $D=1
M467 222 86 440 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=19120 $D=1
M468 441 86 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=14490 $D=1
M469 442 86 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=19120 $D=1
M470 6 87 443 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=14490 $D=1
M471 7 87 444 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=19120 $D=1
M472 445 88 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=14490 $D=1
M473 446 88 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=19120 $D=1
M474 447 87 207 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=14490 $D=1
M475 448 87 208 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=19120 $D=1
M476 6 447 730 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=14490 $D=1
M477 7 448 731 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=19120 $D=1
M478 449 730 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=14490 $D=1
M479 450 731 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=19120 $D=1
M480 447 443 449 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=14490 $D=1
M481 448 444 450 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=19120 $D=1
M482 449 88 217 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=14490 $D=1
M483 450 88 218 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=19120 $D=1
M484 221 89 449 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=14490 $D=1
M485 222 89 450 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=19120 $D=1
M486 451 89 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=14490 $D=1
M487 452 89 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=19120 $D=1
M488 6 90 453 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=14490 $D=1
M489 7 90 454 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=19120 $D=1
M490 455 91 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=14490 $D=1
M491 456 91 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=19120 $D=1
M492 457 90 207 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=14490 $D=1
M493 458 90 208 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=19120 $D=1
M494 6 457 732 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=14490 $D=1
M495 7 458 733 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=19120 $D=1
M496 459 732 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=14490 $D=1
M497 460 733 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=19120 $D=1
M498 457 453 459 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=14490 $D=1
M499 458 454 460 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=19120 $D=1
M500 459 91 217 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=14490 $D=1
M501 460 91 218 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=19120 $D=1
M502 221 92 459 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=14490 $D=1
M503 222 92 460 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=19120 $D=1
M504 461 92 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=14490 $D=1
M505 462 92 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=19120 $D=1
M506 6 93 463 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=14490 $D=1
M507 7 93 464 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=19120 $D=1
M508 465 94 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=14490 $D=1
M509 466 94 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=19120 $D=1
M510 467 93 207 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=14490 $D=1
M511 468 93 208 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=19120 $D=1
M512 6 467 734 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=14490 $D=1
M513 7 468 735 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=19120 $D=1
M514 469 734 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=14490 $D=1
M515 470 735 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=19120 $D=1
M516 467 463 469 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=14490 $D=1
M517 468 464 470 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=19120 $D=1
M518 469 94 217 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=14490 $D=1
M519 470 94 218 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=19120 $D=1
M520 221 95 469 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=14490 $D=1
M521 222 95 470 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=19120 $D=1
M522 471 95 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=14490 $D=1
M523 472 95 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=19120 $D=1
M524 6 96 473 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=14490 $D=1
M525 7 96 474 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=19120 $D=1
M526 475 97 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=14490 $D=1
M527 476 97 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=19120 $D=1
M528 477 96 207 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=14490 $D=1
M529 478 96 208 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=19120 $D=1
M530 6 477 736 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=14490 $D=1
M531 7 478 737 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=19120 $D=1
M532 479 736 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=14490 $D=1
M533 480 737 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=19120 $D=1
M534 477 473 479 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=14490 $D=1
M535 478 474 480 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=19120 $D=1
M536 479 97 217 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=14490 $D=1
M537 480 97 218 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=19120 $D=1
M538 221 98 479 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=14490 $D=1
M539 222 98 480 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=19120 $D=1
M540 481 98 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=14490 $D=1
M541 482 98 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=19120 $D=1
M542 6 99 483 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=14490 $D=1
M543 7 99 484 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=19120 $D=1
M544 485 100 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=14490 $D=1
M545 486 100 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=19120 $D=1
M546 487 99 207 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=14490 $D=1
M547 488 99 208 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=19120 $D=1
M548 6 487 738 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=14490 $D=1
M549 7 488 739 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=19120 $D=1
M550 489 738 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=14490 $D=1
M551 490 739 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=19120 $D=1
M552 487 483 489 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=14490 $D=1
M553 488 484 490 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=19120 $D=1
M554 489 100 217 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=14490 $D=1
M555 490 100 218 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=19120 $D=1
M556 221 101 489 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=14490 $D=1
M557 222 101 490 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=19120 $D=1
M558 491 101 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=14490 $D=1
M559 492 101 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=19120 $D=1
M560 6 102 493 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=14490 $D=1
M561 7 102 494 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=19120 $D=1
M562 495 103 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=14490 $D=1
M563 496 103 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=19120 $D=1
M564 497 102 207 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=14490 $D=1
M565 498 102 208 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=19120 $D=1
M566 6 497 740 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=14490 $D=1
M567 7 498 741 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=19120 $D=1
M568 499 740 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=14490 $D=1
M569 500 741 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=19120 $D=1
M570 497 493 499 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=14490 $D=1
M571 498 494 500 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=19120 $D=1
M572 499 103 217 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=14490 $D=1
M573 500 103 218 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=19120 $D=1
M574 221 104 499 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=14490 $D=1
M575 222 104 500 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=19120 $D=1
M576 501 104 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=14490 $D=1
M577 502 104 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=19120 $D=1
M578 6 105 503 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=14490 $D=1
M579 7 105 504 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=19120 $D=1
M580 505 106 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=14490 $D=1
M581 506 106 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=19120 $D=1
M582 507 105 207 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=14490 $D=1
M583 508 105 208 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=19120 $D=1
M584 6 507 742 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=14490 $D=1
M585 7 508 743 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=19120 $D=1
M586 509 742 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=14490 $D=1
M587 510 743 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=19120 $D=1
M588 507 503 509 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=14490 $D=1
M589 508 504 510 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=19120 $D=1
M590 509 106 217 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=14490 $D=1
M591 510 106 218 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=19120 $D=1
M592 221 107 509 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=14490 $D=1
M593 222 107 510 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=19120 $D=1
M594 511 107 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=14490 $D=1
M595 512 107 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=19120 $D=1
M596 6 108 513 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=14490 $D=1
M597 7 108 514 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=19120 $D=1
M598 515 109 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=14490 $D=1
M599 516 109 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=19120 $D=1
M600 517 108 207 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=14490 $D=1
M601 518 108 208 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=19120 $D=1
M602 6 517 744 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=14490 $D=1
M603 7 518 745 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=19120 $D=1
M604 519 744 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=14490 $D=1
M605 520 745 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=19120 $D=1
M606 517 513 519 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=14490 $D=1
M607 518 514 520 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=19120 $D=1
M608 519 109 217 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=14490 $D=1
M609 520 109 218 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=19120 $D=1
M610 221 110 519 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=14490 $D=1
M611 222 110 520 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=19120 $D=1
M612 521 110 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=14490 $D=1
M613 522 110 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=19120 $D=1
M614 6 111 523 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=14490 $D=1
M615 7 111 524 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=19120 $D=1
M616 525 112 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=14490 $D=1
M617 526 112 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=19120 $D=1
M618 6 112 217 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=14490 $D=1
M619 7 112 218 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=19120 $D=1
M620 221 111 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=14490 $D=1
M621 222 111 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=19120 $D=1
M622 6 529 527 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=14490 $D=1
M623 7 530 528 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=19120 $D=1
M624 529 113 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=14490 $D=1
M625 530 113 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=19120 $D=1
M626 746 217 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=14490 $D=1
M627 747 218 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=19120 $D=1
M628 531 527 746 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=14490 $D=1
M629 532 528 747 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=19120 $D=1
M630 6 531 533 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=14490 $D=1
M631 7 532 534 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=19120 $D=1
M632 748 533 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=14490 $D=1
M633 749 534 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=19120 $D=1
M634 531 529 748 6 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=14490 $D=1
M635 532 530 749 7 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=19120 $D=1
M636 6 537 535 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=14490 $D=1
M637 7 538 536 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=19120 $D=1
M638 537 113 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=14490 $D=1
M639 538 113 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=19120 $D=1
M640 750 221 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=14490 $D=1
M641 751 222 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=19120 $D=1
M642 539 535 750 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=14490 $D=1
M643 540 536 751 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=19120 $D=1
M644 6 539 114 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=14490 $D=1
M645 7 540 115 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=19120 $D=1
M646 752 114 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=14490 $D=1
M647 753 115 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=19120 $D=1
M648 539 537 752 6 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=14490 $D=1
M649 540 538 753 7 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=19120 $D=1
M650 541 116 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=14490 $D=1
M651 542 116 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=19120 $D=1
M652 543 541 533 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=14490 $D=1
M653 544 542 534 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=19120 $D=1
M654 117 116 543 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=14490 $D=1
M655 118 116 544 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=19120 $D=1
M656 545 119 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=14490 $D=1
M657 546 119 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=19120 $D=1
M658 548 545 547 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=14490 $D=1
M659 549 546 115 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=19120 $D=1
M660 754 119 548 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=14490 $D=1
M661 755 119 549 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=19120 $D=1
M662 6 547 754 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=14490 $D=1
M663 7 115 755 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=19120 $D=1
M664 550 120 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=14490 $D=1
M665 551 120 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=19120 $D=1
M666 552 550 548 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=14490 $D=1
M667 553 551 549 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=19120 $D=1
M668 12 120 552 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=14490 $D=1
M669 13 120 553 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=19120 $D=1
M670 555 554 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=14490 $D=1
M671 556 121 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=19120 $D=1
M672 6 559 557 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=14490 $D=1
M673 7 560 558 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=19120 $D=1
M674 561 543 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=14490 $D=1
M675 562 544 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=19120 $D=1
M676 559 561 554 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=14490 $D=1
M677 560 562 121 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=19120 $D=1
M678 555 543 559 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=14490 $D=1
M679 556 544 560 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=19120 $D=1
M680 563 557 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=14490 $D=1
M681 564 558 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=19120 $D=1
M682 122 563 552 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=14490 $D=1
M683 554 564 553 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=19120 $D=1
M684 543 557 122 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=14490 $D=1
M685 544 558 554 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=19120 $D=1
M686 565 122 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=14490 $D=1
M687 566 554 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=19120 $D=1
M688 567 557 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=14490 $D=1
M689 568 558 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=19120 $D=1
M690 569 567 565 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=14490 $D=1
M691 570 568 566 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=19120 $D=1
M692 552 557 569 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=14490 $D=1
M693 553 558 570 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=19120 $D=1
M694 571 543 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=14490 $D=1
M695 572 544 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=19120 $D=1
M696 6 552 571 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=14490 $D=1
M697 7 553 572 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=19120 $D=1
M698 573 569 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=14490 $D=1
M699 574 570 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=19120 $D=1
M700 782 543 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=14490 $D=1
M701 783 544 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=19120 $D=1
M702 575 552 782 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=14490 $D=1
M703 576 553 783 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=19120 $D=1
M704 784 543 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=14490 $D=1
M705 785 544 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=19120 $D=1
M706 577 552 784 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=14490 $D=1
M707 578 553 785 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=19120 $D=1
M708 581 543 579 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=14490 $D=1
M709 582 544 580 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=19120 $D=1
M710 579 552 581 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=14490 $D=1
M711 580 553 582 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=19120 $D=1
M712 6 577 579 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=14490 $D=1
M713 7 578 580 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=19120 $D=1
M714 583 127 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=14490 $D=1
M715 584 127 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=19120 $D=1
M716 585 583 571 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=14490 $D=1
M717 586 584 572 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=19120 $D=1
M718 575 127 585 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=14490 $D=1
M719 576 127 586 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=19120 $D=1
M720 587 583 573 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=14490 $D=1
M721 588 584 574 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=19120 $D=1
M722 581 127 587 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=14490 $D=1
M723 582 127 588 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=19120 $D=1
M724 589 128 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=14490 $D=1
M725 590 128 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=19120 $D=1
M726 591 589 587 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=14490 $D=1
M727 592 590 588 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=19120 $D=1
M728 585 128 591 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=14490 $D=1
M729 586 128 592 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=19120 $D=1
M730 14 591 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=14490 $D=1
M731 15 592 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=19120 $D=1
M732 593 129 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=14490 $D=1
M733 594 129 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=19120 $D=1
M734 595 593 130 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=14490 $D=1
M735 596 594 131 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=19120 $D=1
M736 132 129 595 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=14490 $D=1
M737 133 129 596 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=19120 $D=1
M738 597 129 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=14490 $D=1
M739 598 129 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=19120 $D=1
M740 600 597 134 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=14490 $D=1
M741 601 598 136 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=19120 $D=1
M742 137 129 600 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=14490 $D=1
M743 135 129 601 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=19120 $D=1
M744 602 129 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=14490 $D=1
M745 603 129 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=19120 $D=1
M746 604 602 123 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=14490 $D=1
M747 605 603 126 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=19120 $D=1
M748 138 129 604 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=14490 $D=1
M749 139 129 605 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=19120 $D=1
M750 606 129 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=14490 $D=1
M751 607 129 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=19120 $D=1
M752 608 606 140 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=14490 $D=1
M753 609 607 141 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=19120 $D=1
M754 138 129 608 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=14490 $D=1
M755 138 129 609 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=19120 $D=1
M756 610 129 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=14490 $D=1
M757 611 129 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=19120 $D=1
M758 612 610 142 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=14490 $D=1
M759 613 611 143 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=19120 $D=1
M760 138 129 612 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=14490 $D=1
M761 138 129 613 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=19120 $D=1
M762 6 543 764 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=14490 $D=1
M763 7 544 765 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=19120 $D=1
M764 133 764 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=14490 $D=1
M765 130 765 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=19120 $D=1
M766 614 144 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=14490 $D=1
M767 615 144 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=19120 $D=1
M768 145 614 133 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=14490 $D=1
M769 146 615 130 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=19120 $D=1
M770 595 144 145 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=14490 $D=1
M771 596 144 146 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=19120 $D=1
M772 616 147 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=14490 $D=1
M773 617 147 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=19120 $D=1
M774 148 616 145 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=14490 $D=1
M775 125 617 146 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=19120 $D=1
M776 600 147 148 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=14490 $D=1
M777 601 147 125 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=19120 $D=1
M778 618 149 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=14490 $D=1
M779 619 149 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=19120 $D=1
M780 150 618 148 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=14490 $D=1
M781 151 619 125 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=19120 $D=1
M782 604 149 150 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=14490 $D=1
M783 605 149 151 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=19120 $D=1
M784 620 152 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=14490 $D=1
M785 621 152 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=19120 $D=1
M786 153 620 150 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=14490 $D=1
M787 154 621 151 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=19120 $D=1
M788 608 152 153 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=14490 $D=1
M789 609 152 154 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=19120 $D=1
M790 622 155 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=14490 $D=1
M791 623 155 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=19120 $D=1
M792 193 622 153 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=14490 $D=1
M793 194 623 154 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=19120 $D=1
M794 612 155 193 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=14490 $D=1
M795 613 155 194 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=19120 $D=1
M796 624 156 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=14490 $D=1
M797 625 156 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=19120 $D=1
M798 626 624 547 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=14490 $D=1
M799 627 625 115 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=19120 $D=1
M800 12 156 626 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=14490 $D=1
M801 13 156 627 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=19120 $D=1
M802 786 533 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=14490 $D=1
M803 787 534 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=19120 $D=1
M804 628 626 786 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=14490 $D=1
M805 629 627 787 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=19120 $D=1
M806 632 533 630 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=14490 $D=1
M807 633 534 631 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=19120 $D=1
M808 630 626 632 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=14490 $D=1
M809 631 627 633 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=19120 $D=1
M810 6 628 630 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=14490 $D=1
M811 7 629 631 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=19120 $D=1
M812 788 157 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=14490 $D=1
M813 789 634 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=19120 $D=1
M814 766 632 788 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=14490 $D=1
M815 767 633 789 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=19120 $D=1
M816 634 766 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=14490 $D=1
M817 635 767 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=19120 $D=1
M818 636 533 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=14490 $D=1
M819 637 534 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=19120 $D=1
M820 6 638 636 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=14490 $D=1
M821 7 639 637 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=19120 $D=1
M822 638 626 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=14490 $D=1
M823 639 627 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=19120 $D=1
M824 790 636 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=14490 $D=1
M825 791 637 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=19120 $D=1
M826 640 157 790 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=14490 $D=1
M827 641 634 791 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=19120 $D=1
M828 643 158 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=14490 $D=1
M829 644 642 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=19120 $D=1
M830 792 640 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=14490 $D=1
M831 793 641 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=19120 $D=1
M832 642 643 792 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=14490 $D=1
M833 159 644 793 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=19120 $D=1
M834 646 645 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=14490 $D=1
M835 647 160 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=19120 $D=1
M836 6 650 648 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=14490 $D=1
M837 7 651 649 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=19120 $D=1
M838 652 117 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=14490 $D=1
M839 653 118 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=19120 $D=1
M840 650 652 645 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=14490 $D=1
M841 651 653 160 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=19120 $D=1
M842 646 117 650 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=14490 $D=1
M843 647 118 651 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=19120 $D=1
M844 654 648 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=14490 $D=1
M845 655 649 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=19120 $D=1
M846 161 654 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=14490 $D=1
M847 645 655 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=19120 $D=1
M848 117 648 161 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=14490 $D=1
M849 118 649 645 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=19120 $D=1
M850 656 161 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=14490 $D=1
M851 657 645 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=19120 $D=1
M852 658 648 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=14490 $D=1
M853 659 649 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=19120 $D=1
M854 195 658 656 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=14490 $D=1
M855 196 659 657 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=19120 $D=1
M856 6 648 195 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=14490 $D=1
M857 7 649 196 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=19120 $D=1
M858 660 162 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=14490 $D=1
M859 661 162 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=19120 $D=1
M860 662 660 195 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=14490 $D=1
M861 663 661 196 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=19120 $D=1
M862 14 162 662 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=14490 $D=1
M863 15 162 663 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=19120 $D=1
M864 664 163 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=14490 $D=1
M865 665 163 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=19120 $D=1
M866 163 664 662 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=14490 $D=1
M867 163 665 663 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=19120 $D=1
M868 6 163 163 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=14490 $D=1
M869 7 163 163 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=19120 $D=1
M870 666 113 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=14490 $D=1
M871 667 113 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=19120 $D=1
M872 6 666 668 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=14490 $D=1
M873 7 667 669 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=19120 $D=1
M874 670 113 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=14490 $D=1
M875 671 113 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=19120 $D=1
M876 672 666 163 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=14490 $D=1
M877 673 667 163 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=19120 $D=1
M878 6 672 768 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=14490 $D=1
M879 7 673 769 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=19120 $D=1
M880 674 768 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=14490 $D=1
M881 675 769 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=19120 $D=1
M882 672 668 674 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=14490 $D=1
M883 673 669 675 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=19120 $D=1
M884 676 113 674 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=14490 $D=1
M885 677 113 675 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=19120 $D=1
M886 6 680 678 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=14490 $D=1
M887 7 681 679 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=19120 $D=1
M888 680 113 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=14490 $D=1
M889 681 113 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=19120 $D=1
M890 770 676 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=14490 $D=1
M891 771 677 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=19120 $D=1
M892 682 678 770 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=14490 $D=1
M893 683 679 771 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=19120 $D=1
M894 6 682 117 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=14490 $D=1
M895 7 683 118 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=19120 $D=1
M896 772 117 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=14490 $D=1
M897 773 118 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=19120 $D=1
M898 682 680 772 6 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=14490 $D=1
M899 683 681 773 7 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=19120 $D=1
M900 169 1 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=15740 $D=0
M901 170 1 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=20370 $D=0
M902 171 1 2 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=15740 $D=0
M903 172 1 3 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=20370 $D=0
M904 6 169 171 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=15740 $D=0
M905 7 170 172 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=20370 $D=0
M906 173 1 4 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=15740 $D=0
M907 174 1 4 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=20370 $D=0
M908 5 169 173 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=15740 $D=0
M909 5 170 174 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=20370 $D=0
M910 175 1 6 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=15740 $D=0
M911 176 1 7 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=20370 $D=0
M912 6 169 175 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=15740 $D=0
M913 7 170 176 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=20370 $D=0
M914 179 9 175 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=15740 $D=0
M915 180 9 176 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=20370 $D=0
M916 177 9 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=15740 $D=0
M917 178 9 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=20370 $D=0
M918 181 9 173 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=15740 $D=0
M919 182 9 174 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=20370 $D=0
M920 171 177 181 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=15740 $D=0
M921 172 178 182 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=20370 $D=0
M922 183 10 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=15740 $D=0
M923 184 10 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=20370 $D=0
M924 185 10 181 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=15740 $D=0
M925 186 10 182 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=20370 $D=0
M926 179 183 185 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=15740 $D=0
M927 180 184 186 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=20370 $D=0
M928 187 11 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=15740 $D=0
M929 188 11 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=20370 $D=0
M930 189 11 6 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=15740 $D=0
M931 190 11 7 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=20370 $D=0
M932 12 187 189 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=15740 $D=0
M933 13 188 190 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=20370 $D=0
M934 191 11 14 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=15740 $D=0
M935 192 11 15 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=20370 $D=0
M936 193 187 191 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=15740 $D=0
M937 194 188 192 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=20370 $D=0
M938 197 11 195 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=15740 $D=0
M939 198 11 196 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=20370 $D=0
M940 185 187 197 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=15740 $D=0
M941 186 188 198 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=20370 $D=0
M942 201 16 197 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=15740 $D=0
M943 202 16 198 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=20370 $D=0
M944 199 16 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=15740 $D=0
M945 200 16 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=20370 $D=0
M946 203 16 191 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=15740 $D=0
M947 204 16 192 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=20370 $D=0
M948 189 199 203 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=15740 $D=0
M949 190 200 204 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=20370 $D=0
M950 205 17 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=15740 $D=0
M951 206 17 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=20370 $D=0
M952 207 17 203 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=15740 $D=0
M953 208 17 204 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=20370 $D=0
M954 201 205 207 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=15740 $D=0
M955 202 206 208 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=20370 $D=0
M956 164 18 209 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=15740 $D=0
M957 165 18 210 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=20370 $D=0
M958 211 19 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=15740 $D=0
M959 212 19 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=20370 $D=0
M960 213 209 207 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=15740 $D=0
M961 214 210 208 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=20370 $D=0
M962 164 213 684 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=15740 $D=0
M963 165 214 685 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=20370 $D=0
M964 215 684 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=15740 $D=0
M965 216 685 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=20370 $D=0
M966 213 18 215 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=15740 $D=0
M967 214 18 216 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=20370 $D=0
M968 215 211 217 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=15740 $D=0
M969 216 212 218 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=20370 $D=0
M970 221 219 215 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=15740 $D=0
M971 222 220 216 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=20370 $D=0
M972 219 20 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=15740 $D=0
M973 220 20 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=20370 $D=0
M974 164 21 223 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=15740 $D=0
M975 165 21 224 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=20370 $D=0
M976 225 22 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=15740 $D=0
M977 226 22 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=20370 $D=0
M978 227 223 207 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=15740 $D=0
M979 228 224 208 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=20370 $D=0
M980 164 227 686 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=15740 $D=0
M981 165 228 687 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=20370 $D=0
M982 229 686 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=15740 $D=0
M983 230 687 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=20370 $D=0
M984 227 21 229 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=15740 $D=0
M985 228 21 230 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=20370 $D=0
M986 229 225 217 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=15740 $D=0
M987 230 226 218 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=20370 $D=0
M988 221 231 229 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=15740 $D=0
M989 222 232 230 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=20370 $D=0
M990 231 23 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=15740 $D=0
M991 232 23 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=20370 $D=0
M992 164 24 233 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=15740 $D=0
M993 165 24 234 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=20370 $D=0
M994 235 25 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=15740 $D=0
M995 236 25 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=20370 $D=0
M996 237 233 207 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=15740 $D=0
M997 238 234 208 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=20370 $D=0
M998 164 237 688 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=15740 $D=0
M999 165 238 689 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=20370 $D=0
M1000 239 688 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=15740 $D=0
M1001 240 689 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=20370 $D=0
M1002 237 24 239 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=15740 $D=0
M1003 238 24 240 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=20370 $D=0
M1004 239 235 217 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=15740 $D=0
M1005 240 236 218 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=20370 $D=0
M1006 221 241 239 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=15740 $D=0
M1007 222 242 240 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=20370 $D=0
M1008 241 26 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=15740 $D=0
M1009 242 26 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=20370 $D=0
M1010 164 27 243 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=15740 $D=0
M1011 165 27 244 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=20370 $D=0
M1012 245 28 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=15740 $D=0
M1013 246 28 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=20370 $D=0
M1014 247 243 207 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=15740 $D=0
M1015 248 244 208 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=20370 $D=0
M1016 164 247 690 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=15740 $D=0
M1017 165 248 691 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=20370 $D=0
M1018 249 690 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=15740 $D=0
M1019 250 691 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=20370 $D=0
M1020 247 27 249 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=15740 $D=0
M1021 248 27 250 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=20370 $D=0
M1022 249 245 217 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=15740 $D=0
M1023 250 246 218 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=20370 $D=0
M1024 221 251 249 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=15740 $D=0
M1025 222 252 250 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=20370 $D=0
M1026 251 29 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=15740 $D=0
M1027 252 29 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=20370 $D=0
M1028 164 30 253 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=15740 $D=0
M1029 165 30 254 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=20370 $D=0
M1030 255 31 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=15740 $D=0
M1031 256 31 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=20370 $D=0
M1032 257 253 207 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=15740 $D=0
M1033 258 254 208 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=20370 $D=0
M1034 164 257 692 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=15740 $D=0
M1035 165 258 693 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=20370 $D=0
M1036 259 692 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=15740 $D=0
M1037 260 693 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=20370 $D=0
M1038 257 30 259 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=15740 $D=0
M1039 258 30 260 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=20370 $D=0
M1040 259 255 217 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=15740 $D=0
M1041 260 256 218 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=20370 $D=0
M1042 221 261 259 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=15740 $D=0
M1043 222 262 260 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=20370 $D=0
M1044 261 32 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=15740 $D=0
M1045 262 32 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=20370 $D=0
M1046 164 33 263 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=15740 $D=0
M1047 165 33 264 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=20370 $D=0
M1048 265 34 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=15740 $D=0
M1049 266 34 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=20370 $D=0
M1050 267 263 207 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=15740 $D=0
M1051 268 264 208 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=20370 $D=0
M1052 164 267 694 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=15740 $D=0
M1053 165 268 695 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=20370 $D=0
M1054 269 694 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=15740 $D=0
M1055 270 695 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=20370 $D=0
M1056 267 33 269 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=15740 $D=0
M1057 268 33 270 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=20370 $D=0
M1058 269 265 217 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=15740 $D=0
M1059 270 266 218 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=20370 $D=0
M1060 221 271 269 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=15740 $D=0
M1061 222 272 270 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=20370 $D=0
M1062 271 35 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=15740 $D=0
M1063 272 35 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=20370 $D=0
M1064 164 36 273 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=15740 $D=0
M1065 165 36 274 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=20370 $D=0
M1066 275 37 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=15740 $D=0
M1067 276 37 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=20370 $D=0
M1068 277 273 207 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=15740 $D=0
M1069 278 274 208 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=20370 $D=0
M1070 164 277 696 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=15740 $D=0
M1071 165 278 697 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=20370 $D=0
M1072 279 696 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=15740 $D=0
M1073 280 697 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=20370 $D=0
M1074 277 36 279 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=15740 $D=0
M1075 278 36 280 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=20370 $D=0
M1076 279 275 217 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=15740 $D=0
M1077 280 276 218 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=20370 $D=0
M1078 221 281 279 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=15740 $D=0
M1079 222 282 280 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=20370 $D=0
M1080 281 38 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=15740 $D=0
M1081 282 38 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=20370 $D=0
M1082 164 39 283 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=15740 $D=0
M1083 165 39 284 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=20370 $D=0
M1084 285 40 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=15740 $D=0
M1085 286 40 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=20370 $D=0
M1086 287 283 207 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=15740 $D=0
M1087 288 284 208 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=20370 $D=0
M1088 164 287 698 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=15740 $D=0
M1089 165 288 699 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=20370 $D=0
M1090 289 698 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=15740 $D=0
M1091 290 699 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=20370 $D=0
M1092 287 39 289 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=15740 $D=0
M1093 288 39 290 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=20370 $D=0
M1094 289 285 217 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=15740 $D=0
M1095 290 286 218 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=20370 $D=0
M1096 221 291 289 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=15740 $D=0
M1097 222 292 290 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=20370 $D=0
M1098 291 41 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=15740 $D=0
M1099 292 41 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=20370 $D=0
M1100 164 42 293 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=15740 $D=0
M1101 165 42 294 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=20370 $D=0
M1102 295 43 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=15740 $D=0
M1103 296 43 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=20370 $D=0
M1104 297 293 207 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=15740 $D=0
M1105 298 294 208 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=20370 $D=0
M1106 164 297 700 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=15740 $D=0
M1107 165 298 701 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=20370 $D=0
M1108 299 700 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=15740 $D=0
M1109 300 701 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=20370 $D=0
M1110 297 42 299 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=15740 $D=0
M1111 298 42 300 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=20370 $D=0
M1112 299 295 217 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=15740 $D=0
M1113 300 296 218 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=20370 $D=0
M1114 221 301 299 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=15740 $D=0
M1115 222 302 300 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=20370 $D=0
M1116 301 44 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=15740 $D=0
M1117 302 44 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=20370 $D=0
M1118 164 45 303 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=15740 $D=0
M1119 165 45 304 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=20370 $D=0
M1120 305 46 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=15740 $D=0
M1121 306 46 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=20370 $D=0
M1122 307 303 207 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=15740 $D=0
M1123 308 304 208 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=20370 $D=0
M1124 164 307 702 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=15740 $D=0
M1125 165 308 703 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=20370 $D=0
M1126 309 702 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=15740 $D=0
M1127 310 703 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=20370 $D=0
M1128 307 45 309 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=15740 $D=0
M1129 308 45 310 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=20370 $D=0
M1130 309 305 217 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=15740 $D=0
M1131 310 306 218 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=20370 $D=0
M1132 221 311 309 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=15740 $D=0
M1133 222 312 310 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=20370 $D=0
M1134 311 47 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=15740 $D=0
M1135 312 47 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=20370 $D=0
M1136 164 48 313 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=15740 $D=0
M1137 165 48 314 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=20370 $D=0
M1138 315 49 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=15740 $D=0
M1139 316 49 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=20370 $D=0
M1140 317 313 207 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=15740 $D=0
M1141 318 314 208 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=20370 $D=0
M1142 164 317 704 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=15740 $D=0
M1143 165 318 705 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=20370 $D=0
M1144 319 704 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=15740 $D=0
M1145 320 705 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=20370 $D=0
M1146 317 48 319 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=15740 $D=0
M1147 318 48 320 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=20370 $D=0
M1148 319 315 217 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=15740 $D=0
M1149 320 316 218 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=20370 $D=0
M1150 221 321 319 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=15740 $D=0
M1151 222 322 320 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=20370 $D=0
M1152 321 50 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=15740 $D=0
M1153 322 50 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=20370 $D=0
M1154 164 51 323 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=15740 $D=0
M1155 165 51 324 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=20370 $D=0
M1156 325 52 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=15740 $D=0
M1157 326 52 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=20370 $D=0
M1158 327 323 207 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=15740 $D=0
M1159 328 324 208 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=20370 $D=0
M1160 164 327 706 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=15740 $D=0
M1161 165 328 707 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=20370 $D=0
M1162 329 706 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=15740 $D=0
M1163 330 707 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=20370 $D=0
M1164 327 51 329 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=15740 $D=0
M1165 328 51 330 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=20370 $D=0
M1166 329 325 217 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=15740 $D=0
M1167 330 326 218 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=20370 $D=0
M1168 221 331 329 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=15740 $D=0
M1169 222 332 330 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=20370 $D=0
M1170 331 53 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=15740 $D=0
M1171 332 53 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=20370 $D=0
M1172 164 54 333 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=15740 $D=0
M1173 165 54 334 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=20370 $D=0
M1174 335 55 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=15740 $D=0
M1175 336 55 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=20370 $D=0
M1176 337 333 207 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=15740 $D=0
M1177 338 334 208 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=20370 $D=0
M1178 164 337 708 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=15740 $D=0
M1179 165 338 709 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=20370 $D=0
M1180 339 708 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=15740 $D=0
M1181 340 709 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=20370 $D=0
M1182 337 54 339 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=15740 $D=0
M1183 338 54 340 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=20370 $D=0
M1184 339 335 217 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=15740 $D=0
M1185 340 336 218 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=20370 $D=0
M1186 221 341 339 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=15740 $D=0
M1187 222 342 340 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=20370 $D=0
M1188 341 56 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=15740 $D=0
M1189 342 56 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=20370 $D=0
M1190 164 57 343 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=15740 $D=0
M1191 165 57 344 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=20370 $D=0
M1192 345 58 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=15740 $D=0
M1193 346 58 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=20370 $D=0
M1194 347 343 207 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=15740 $D=0
M1195 348 344 208 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=20370 $D=0
M1196 164 347 710 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=15740 $D=0
M1197 165 348 711 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=20370 $D=0
M1198 349 710 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=15740 $D=0
M1199 350 711 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=20370 $D=0
M1200 347 57 349 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=15740 $D=0
M1201 348 57 350 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=20370 $D=0
M1202 349 345 217 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=15740 $D=0
M1203 350 346 218 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=20370 $D=0
M1204 221 351 349 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=15740 $D=0
M1205 222 352 350 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=20370 $D=0
M1206 351 59 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=15740 $D=0
M1207 352 59 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=20370 $D=0
M1208 164 60 353 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=15740 $D=0
M1209 165 60 354 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=20370 $D=0
M1210 355 61 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=15740 $D=0
M1211 356 61 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=20370 $D=0
M1212 357 353 207 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=15740 $D=0
M1213 358 354 208 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=20370 $D=0
M1214 164 357 712 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=15740 $D=0
M1215 165 358 713 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=20370 $D=0
M1216 359 712 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=15740 $D=0
M1217 360 713 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=20370 $D=0
M1218 357 60 359 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=15740 $D=0
M1219 358 60 360 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=20370 $D=0
M1220 359 355 217 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=15740 $D=0
M1221 360 356 218 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=20370 $D=0
M1222 221 361 359 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=15740 $D=0
M1223 222 362 360 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=20370 $D=0
M1224 361 62 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=15740 $D=0
M1225 362 62 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=20370 $D=0
M1226 164 63 363 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=15740 $D=0
M1227 165 63 364 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=20370 $D=0
M1228 365 64 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=15740 $D=0
M1229 366 64 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=20370 $D=0
M1230 367 363 207 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=15740 $D=0
M1231 368 364 208 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=20370 $D=0
M1232 164 367 714 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=15740 $D=0
M1233 165 368 715 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=20370 $D=0
M1234 369 714 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=15740 $D=0
M1235 370 715 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=20370 $D=0
M1236 367 63 369 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=15740 $D=0
M1237 368 63 370 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=20370 $D=0
M1238 369 365 217 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=15740 $D=0
M1239 370 366 218 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=20370 $D=0
M1240 221 371 369 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=15740 $D=0
M1241 222 372 370 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=20370 $D=0
M1242 371 65 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=15740 $D=0
M1243 372 65 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=20370 $D=0
M1244 164 66 373 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=15740 $D=0
M1245 165 66 374 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=20370 $D=0
M1246 375 67 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=15740 $D=0
M1247 376 67 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=20370 $D=0
M1248 377 373 207 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=15740 $D=0
M1249 378 374 208 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=20370 $D=0
M1250 164 377 716 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=15740 $D=0
M1251 165 378 717 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=20370 $D=0
M1252 379 716 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=15740 $D=0
M1253 380 717 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=20370 $D=0
M1254 377 66 379 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=15740 $D=0
M1255 378 66 380 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=20370 $D=0
M1256 379 375 217 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=15740 $D=0
M1257 380 376 218 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=20370 $D=0
M1258 221 381 379 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=15740 $D=0
M1259 222 382 380 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=20370 $D=0
M1260 381 68 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=15740 $D=0
M1261 382 68 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=20370 $D=0
M1262 164 69 383 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=15740 $D=0
M1263 165 69 384 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=20370 $D=0
M1264 385 70 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=15740 $D=0
M1265 386 70 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=20370 $D=0
M1266 387 383 207 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=15740 $D=0
M1267 388 384 208 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=20370 $D=0
M1268 164 387 718 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=15740 $D=0
M1269 165 388 719 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=20370 $D=0
M1270 389 718 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=15740 $D=0
M1271 390 719 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=20370 $D=0
M1272 387 69 389 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=15740 $D=0
M1273 388 69 390 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=20370 $D=0
M1274 389 385 217 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=15740 $D=0
M1275 390 386 218 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=20370 $D=0
M1276 221 391 389 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=15740 $D=0
M1277 222 392 390 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=20370 $D=0
M1278 391 71 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=15740 $D=0
M1279 392 71 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=20370 $D=0
M1280 164 72 393 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=15740 $D=0
M1281 165 72 394 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=20370 $D=0
M1282 395 73 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=15740 $D=0
M1283 396 73 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=20370 $D=0
M1284 397 393 207 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=15740 $D=0
M1285 398 394 208 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=20370 $D=0
M1286 164 397 720 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=15740 $D=0
M1287 165 398 721 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=20370 $D=0
M1288 399 720 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=15740 $D=0
M1289 400 721 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=20370 $D=0
M1290 397 72 399 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=15740 $D=0
M1291 398 72 400 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=20370 $D=0
M1292 399 395 217 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=15740 $D=0
M1293 400 396 218 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=20370 $D=0
M1294 221 401 399 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=15740 $D=0
M1295 222 402 400 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=20370 $D=0
M1296 401 74 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=15740 $D=0
M1297 402 74 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=20370 $D=0
M1298 164 75 403 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=15740 $D=0
M1299 165 75 404 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=20370 $D=0
M1300 405 76 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=15740 $D=0
M1301 406 76 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=20370 $D=0
M1302 407 403 207 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=15740 $D=0
M1303 408 404 208 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=20370 $D=0
M1304 164 407 722 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=15740 $D=0
M1305 165 408 723 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=20370 $D=0
M1306 409 722 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=15740 $D=0
M1307 410 723 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=20370 $D=0
M1308 407 75 409 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=15740 $D=0
M1309 408 75 410 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=20370 $D=0
M1310 409 405 217 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=15740 $D=0
M1311 410 406 218 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=20370 $D=0
M1312 221 411 409 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=15740 $D=0
M1313 222 412 410 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=20370 $D=0
M1314 411 77 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=15740 $D=0
M1315 412 77 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=20370 $D=0
M1316 164 78 413 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=15740 $D=0
M1317 165 78 414 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=20370 $D=0
M1318 415 79 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=15740 $D=0
M1319 416 79 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=20370 $D=0
M1320 417 413 207 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=15740 $D=0
M1321 418 414 208 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=20370 $D=0
M1322 164 417 724 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=15740 $D=0
M1323 165 418 725 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=20370 $D=0
M1324 419 724 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=15740 $D=0
M1325 420 725 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=20370 $D=0
M1326 417 78 419 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=15740 $D=0
M1327 418 78 420 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=20370 $D=0
M1328 419 415 217 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=15740 $D=0
M1329 420 416 218 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=20370 $D=0
M1330 221 421 419 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=15740 $D=0
M1331 222 422 420 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=20370 $D=0
M1332 421 80 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=15740 $D=0
M1333 422 80 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=20370 $D=0
M1334 164 81 423 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=15740 $D=0
M1335 165 81 424 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=20370 $D=0
M1336 425 82 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=15740 $D=0
M1337 426 82 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=20370 $D=0
M1338 427 423 207 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=15740 $D=0
M1339 428 424 208 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=20370 $D=0
M1340 164 427 726 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=15740 $D=0
M1341 165 428 727 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=20370 $D=0
M1342 429 726 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=15740 $D=0
M1343 430 727 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=20370 $D=0
M1344 427 81 429 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=15740 $D=0
M1345 428 81 430 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=20370 $D=0
M1346 429 425 217 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=15740 $D=0
M1347 430 426 218 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=20370 $D=0
M1348 221 431 429 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=15740 $D=0
M1349 222 432 430 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=20370 $D=0
M1350 431 83 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=15740 $D=0
M1351 432 83 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=20370 $D=0
M1352 164 84 433 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=15740 $D=0
M1353 165 84 434 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=20370 $D=0
M1354 435 85 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=15740 $D=0
M1355 436 85 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=20370 $D=0
M1356 437 433 207 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=15740 $D=0
M1357 438 434 208 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=20370 $D=0
M1358 164 437 728 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=15740 $D=0
M1359 165 438 729 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=20370 $D=0
M1360 439 728 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=15740 $D=0
M1361 440 729 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=20370 $D=0
M1362 437 84 439 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=15740 $D=0
M1363 438 84 440 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=20370 $D=0
M1364 439 435 217 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=15740 $D=0
M1365 440 436 218 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=20370 $D=0
M1366 221 441 439 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=15740 $D=0
M1367 222 442 440 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=20370 $D=0
M1368 441 86 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=15740 $D=0
M1369 442 86 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=20370 $D=0
M1370 164 87 443 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=15740 $D=0
M1371 165 87 444 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=20370 $D=0
M1372 445 88 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=15740 $D=0
M1373 446 88 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=20370 $D=0
M1374 447 443 207 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=15740 $D=0
M1375 448 444 208 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=20370 $D=0
M1376 164 447 730 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=15740 $D=0
M1377 165 448 731 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=20370 $D=0
M1378 449 730 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=15740 $D=0
M1379 450 731 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=20370 $D=0
M1380 447 87 449 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=15740 $D=0
M1381 448 87 450 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=20370 $D=0
M1382 449 445 217 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=15740 $D=0
M1383 450 446 218 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=20370 $D=0
M1384 221 451 449 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=15740 $D=0
M1385 222 452 450 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=20370 $D=0
M1386 451 89 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=15740 $D=0
M1387 452 89 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=20370 $D=0
M1388 164 90 453 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=15740 $D=0
M1389 165 90 454 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=20370 $D=0
M1390 455 91 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=15740 $D=0
M1391 456 91 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=20370 $D=0
M1392 457 453 207 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=15740 $D=0
M1393 458 454 208 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=20370 $D=0
M1394 164 457 732 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=15740 $D=0
M1395 165 458 733 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=20370 $D=0
M1396 459 732 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=15740 $D=0
M1397 460 733 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=20370 $D=0
M1398 457 90 459 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=15740 $D=0
M1399 458 90 460 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=20370 $D=0
M1400 459 455 217 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=15740 $D=0
M1401 460 456 218 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=20370 $D=0
M1402 221 461 459 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=15740 $D=0
M1403 222 462 460 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=20370 $D=0
M1404 461 92 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=15740 $D=0
M1405 462 92 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=20370 $D=0
M1406 164 93 463 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=15740 $D=0
M1407 165 93 464 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=20370 $D=0
M1408 465 94 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=15740 $D=0
M1409 466 94 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=20370 $D=0
M1410 467 463 207 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=15740 $D=0
M1411 468 464 208 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=20370 $D=0
M1412 164 467 734 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=15740 $D=0
M1413 165 468 735 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=20370 $D=0
M1414 469 734 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=15740 $D=0
M1415 470 735 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=20370 $D=0
M1416 467 93 469 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=15740 $D=0
M1417 468 93 470 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=20370 $D=0
M1418 469 465 217 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=15740 $D=0
M1419 470 466 218 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=20370 $D=0
M1420 221 471 469 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=15740 $D=0
M1421 222 472 470 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=20370 $D=0
M1422 471 95 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=15740 $D=0
M1423 472 95 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=20370 $D=0
M1424 164 96 473 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=15740 $D=0
M1425 165 96 474 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=20370 $D=0
M1426 475 97 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=15740 $D=0
M1427 476 97 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=20370 $D=0
M1428 477 473 207 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=15740 $D=0
M1429 478 474 208 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=20370 $D=0
M1430 164 477 736 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=15740 $D=0
M1431 165 478 737 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=20370 $D=0
M1432 479 736 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=15740 $D=0
M1433 480 737 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=20370 $D=0
M1434 477 96 479 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=15740 $D=0
M1435 478 96 480 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=20370 $D=0
M1436 479 475 217 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=15740 $D=0
M1437 480 476 218 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=20370 $D=0
M1438 221 481 479 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=15740 $D=0
M1439 222 482 480 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=20370 $D=0
M1440 481 98 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=15740 $D=0
M1441 482 98 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=20370 $D=0
M1442 164 99 483 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=15740 $D=0
M1443 165 99 484 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=20370 $D=0
M1444 485 100 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=15740 $D=0
M1445 486 100 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=20370 $D=0
M1446 487 483 207 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=15740 $D=0
M1447 488 484 208 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=20370 $D=0
M1448 164 487 738 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=15740 $D=0
M1449 165 488 739 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=20370 $D=0
M1450 489 738 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=15740 $D=0
M1451 490 739 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=20370 $D=0
M1452 487 99 489 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=15740 $D=0
M1453 488 99 490 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=20370 $D=0
M1454 489 485 217 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=15740 $D=0
M1455 490 486 218 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=20370 $D=0
M1456 221 491 489 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=15740 $D=0
M1457 222 492 490 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=20370 $D=0
M1458 491 101 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=15740 $D=0
M1459 492 101 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=20370 $D=0
M1460 164 102 493 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=15740 $D=0
M1461 165 102 494 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=20370 $D=0
M1462 495 103 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=15740 $D=0
M1463 496 103 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=20370 $D=0
M1464 497 493 207 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=15740 $D=0
M1465 498 494 208 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=20370 $D=0
M1466 164 497 740 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=15740 $D=0
M1467 165 498 741 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=20370 $D=0
M1468 499 740 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=15740 $D=0
M1469 500 741 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=20370 $D=0
M1470 497 102 499 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=15740 $D=0
M1471 498 102 500 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=20370 $D=0
M1472 499 495 217 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=15740 $D=0
M1473 500 496 218 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=20370 $D=0
M1474 221 501 499 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=15740 $D=0
M1475 222 502 500 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=20370 $D=0
M1476 501 104 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=15740 $D=0
M1477 502 104 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=20370 $D=0
M1478 164 105 503 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=15740 $D=0
M1479 165 105 504 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=20370 $D=0
M1480 505 106 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=15740 $D=0
M1481 506 106 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=20370 $D=0
M1482 507 503 207 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=15740 $D=0
M1483 508 504 208 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=20370 $D=0
M1484 164 507 742 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=15740 $D=0
M1485 165 508 743 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=20370 $D=0
M1486 509 742 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=15740 $D=0
M1487 510 743 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=20370 $D=0
M1488 507 105 509 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=15740 $D=0
M1489 508 105 510 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=20370 $D=0
M1490 509 505 217 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=15740 $D=0
M1491 510 506 218 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=20370 $D=0
M1492 221 511 509 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=15740 $D=0
M1493 222 512 510 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=20370 $D=0
M1494 511 107 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=15740 $D=0
M1495 512 107 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=20370 $D=0
M1496 164 108 513 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=15740 $D=0
M1497 165 108 514 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=20370 $D=0
M1498 515 109 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=15740 $D=0
M1499 516 109 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=20370 $D=0
M1500 517 513 207 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=15740 $D=0
M1501 518 514 208 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=20370 $D=0
M1502 164 517 744 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=15740 $D=0
M1503 165 518 745 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=20370 $D=0
M1504 519 744 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=15740 $D=0
M1505 520 745 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=20370 $D=0
M1506 517 108 519 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=15740 $D=0
M1507 518 108 520 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=20370 $D=0
M1508 519 515 217 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=15740 $D=0
M1509 520 516 218 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=20370 $D=0
M1510 221 521 519 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=15740 $D=0
M1511 222 522 520 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=20370 $D=0
M1512 521 110 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=15740 $D=0
M1513 522 110 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=20370 $D=0
M1514 164 111 523 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=15740 $D=0
M1515 165 111 524 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=20370 $D=0
M1516 525 112 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=15740 $D=0
M1517 526 112 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=20370 $D=0
M1518 6 525 217 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=15740 $D=0
M1519 7 526 218 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=20370 $D=0
M1520 221 523 6 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=15740 $D=0
M1521 222 524 7 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=20370 $D=0
M1522 164 529 527 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=15740 $D=0
M1523 165 530 528 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=20370 $D=0
M1524 529 113 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=15740 $D=0
M1525 530 113 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=20370 $D=0
M1526 746 217 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=15740 $D=0
M1527 747 218 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=20370 $D=0
M1528 531 529 746 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=15740 $D=0
M1529 532 530 747 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=20370 $D=0
M1530 164 531 533 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=15740 $D=0
M1531 165 532 534 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=20370 $D=0
M1532 748 533 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=15740 $D=0
M1533 749 534 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=20370 $D=0
M1534 531 527 748 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=15740 $D=0
M1535 532 528 749 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=20370 $D=0
M1536 164 537 535 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=15740 $D=0
M1537 165 538 536 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=20370 $D=0
M1538 537 113 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=15740 $D=0
M1539 538 113 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=20370 $D=0
M1540 750 221 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=15740 $D=0
M1541 751 222 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=20370 $D=0
M1542 539 537 750 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=15740 $D=0
M1543 540 538 751 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=20370 $D=0
M1544 164 539 114 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=15740 $D=0
M1545 165 540 115 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=20370 $D=0
M1546 752 114 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=15740 $D=0
M1547 753 115 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=20370 $D=0
M1548 539 535 752 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=15740 $D=0
M1549 540 536 753 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=20370 $D=0
M1550 541 116 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=15740 $D=0
M1551 542 116 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=20370 $D=0
M1552 543 116 533 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=15740 $D=0
M1553 544 116 534 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=20370 $D=0
M1554 117 541 543 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=15740 $D=0
M1555 118 542 544 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=20370 $D=0
M1556 545 119 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=15740 $D=0
M1557 546 119 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=20370 $D=0
M1558 548 119 547 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=15740 $D=0
M1559 549 119 115 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=20370 $D=0
M1560 754 545 548 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=15740 $D=0
M1561 755 546 549 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=20370 $D=0
M1562 164 547 754 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=15740 $D=0
M1563 165 115 755 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=20370 $D=0
M1564 550 120 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=15740 $D=0
M1565 551 120 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=20370 $D=0
M1566 552 120 548 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=15740 $D=0
M1567 553 120 549 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=20370 $D=0
M1568 12 550 552 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=15740 $D=0
M1569 13 551 553 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=20370 $D=0
M1570 555 554 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=15740 $D=0
M1571 556 121 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=20370 $D=0
M1572 164 559 557 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=15740 $D=0
M1573 165 560 558 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=20370 $D=0
M1574 561 543 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=15740 $D=0
M1575 562 544 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=20370 $D=0
M1576 559 543 554 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=15740 $D=0
M1577 560 544 121 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=20370 $D=0
M1578 555 561 559 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=15740 $D=0
M1579 556 562 560 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=20370 $D=0
M1580 563 557 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=15740 $D=0
M1581 564 558 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=20370 $D=0
M1582 122 557 552 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=15740 $D=0
M1583 554 558 553 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=20370 $D=0
M1584 543 563 122 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=15740 $D=0
M1585 544 564 554 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=20370 $D=0
M1586 565 122 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=15740 $D=0
M1587 566 554 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=20370 $D=0
M1588 567 557 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=15740 $D=0
M1589 568 558 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=20370 $D=0
M1590 569 557 565 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=15740 $D=0
M1591 570 558 566 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=20370 $D=0
M1592 552 567 569 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=15740 $D=0
M1593 553 568 570 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=20370 $D=0
M1594 774 543 164 164 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=15380 $D=0
M1595 775 544 165 165 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=20010 $D=0
M1596 571 552 774 164 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=15380 $D=0
M1597 572 553 775 165 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=20010 $D=0
M1598 573 569 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=15740 $D=0
M1599 574 570 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=20370 $D=0
M1600 575 543 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=15740 $D=0
M1601 576 544 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=20370 $D=0
M1602 164 552 575 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=15740 $D=0
M1603 165 553 576 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=20370 $D=0
M1604 577 543 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=15740 $D=0
M1605 578 544 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=20370 $D=0
M1606 164 552 577 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=15740 $D=0
M1607 165 553 578 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=20370 $D=0
M1608 776 543 164 164 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=15560 $D=0
M1609 777 544 165 165 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=20190 $D=0
M1610 581 552 776 164 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=15560 $D=0
M1611 582 553 777 165 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=20190 $D=0
M1612 164 577 581 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=15740 $D=0
M1613 165 578 582 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=20370 $D=0
M1614 583 127 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=15740 $D=0
M1615 584 127 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=20370 $D=0
M1616 585 127 571 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=15740 $D=0
M1617 586 127 572 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=20370 $D=0
M1618 575 583 585 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=15740 $D=0
M1619 576 584 586 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=20370 $D=0
M1620 587 127 573 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=15740 $D=0
M1621 588 127 574 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=20370 $D=0
M1622 581 583 587 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=15740 $D=0
M1623 582 584 588 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=20370 $D=0
M1624 589 128 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=15740 $D=0
M1625 590 128 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=20370 $D=0
M1626 591 128 587 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=15740 $D=0
M1627 592 128 588 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=20370 $D=0
M1628 585 589 591 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=15740 $D=0
M1629 586 590 592 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=20370 $D=0
M1630 14 591 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=15740 $D=0
M1631 15 592 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=20370 $D=0
M1632 593 129 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=15740 $D=0
M1633 594 129 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=20370 $D=0
M1634 595 129 130 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=15740 $D=0
M1635 596 129 131 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=20370 $D=0
M1636 132 593 595 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=15740 $D=0
M1637 133 594 596 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=20370 $D=0
M1638 597 129 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=15740 $D=0
M1639 598 129 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=20370 $D=0
M1640 600 129 134 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=15740 $D=0
M1641 601 129 136 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=20370 $D=0
M1642 137 597 600 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=15740 $D=0
M1643 135 598 601 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=20370 $D=0
M1644 602 129 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=15740 $D=0
M1645 603 129 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=20370 $D=0
M1646 604 129 123 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=15740 $D=0
M1647 605 129 126 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=20370 $D=0
M1648 138 602 604 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=15740 $D=0
M1649 139 603 605 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=20370 $D=0
M1650 606 129 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=15740 $D=0
M1651 607 129 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=20370 $D=0
M1652 608 129 140 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=15740 $D=0
M1653 609 129 141 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=20370 $D=0
M1654 138 606 608 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=15740 $D=0
M1655 138 607 609 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=20370 $D=0
M1656 610 129 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=15740 $D=0
M1657 611 129 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=20370 $D=0
M1658 612 129 142 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=15740 $D=0
M1659 613 129 143 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=20370 $D=0
M1660 138 610 612 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=15740 $D=0
M1661 138 611 613 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=20370 $D=0
M1662 164 543 764 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=15740 $D=0
M1663 165 544 765 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=20370 $D=0
M1664 133 764 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=15740 $D=0
M1665 130 765 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=20370 $D=0
M1666 614 144 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=15740 $D=0
M1667 615 144 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=20370 $D=0
M1668 145 144 133 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=15740 $D=0
M1669 146 144 130 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=20370 $D=0
M1670 595 614 145 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=15740 $D=0
M1671 596 615 146 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=20370 $D=0
M1672 616 147 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=15740 $D=0
M1673 617 147 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=20370 $D=0
M1674 148 147 145 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=15740 $D=0
M1675 125 147 146 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=20370 $D=0
M1676 600 616 148 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=15740 $D=0
M1677 601 617 125 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=20370 $D=0
M1678 618 149 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=15740 $D=0
M1679 619 149 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=20370 $D=0
M1680 150 149 148 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=15740 $D=0
M1681 151 149 125 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=20370 $D=0
M1682 604 618 150 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=15740 $D=0
M1683 605 619 151 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=20370 $D=0
M1684 620 152 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=15740 $D=0
M1685 621 152 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=20370 $D=0
M1686 153 152 150 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=15740 $D=0
M1687 154 152 151 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=20370 $D=0
M1688 608 620 153 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=15740 $D=0
M1689 609 621 154 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=20370 $D=0
M1690 622 155 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=15740 $D=0
M1691 623 155 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=20370 $D=0
M1692 193 155 153 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=15740 $D=0
M1693 194 155 154 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=20370 $D=0
M1694 612 622 193 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=15740 $D=0
M1695 613 623 194 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=20370 $D=0
M1696 624 156 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=15740 $D=0
M1697 625 156 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=20370 $D=0
M1698 626 156 547 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=15740 $D=0
M1699 627 156 115 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=20370 $D=0
M1700 12 624 626 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=15740 $D=0
M1701 13 625 627 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=20370 $D=0
M1702 628 533 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=15740 $D=0
M1703 629 534 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=20370 $D=0
M1704 164 626 628 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=15740 $D=0
M1705 165 627 629 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=20370 $D=0
M1706 778 533 164 164 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=15560 $D=0
M1707 779 534 165 165 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=20190 $D=0
M1708 632 626 778 164 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=15560 $D=0
M1709 633 627 779 165 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=20190 $D=0
M1710 164 628 632 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=15740 $D=0
M1711 165 629 633 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=20370 $D=0
M1712 766 157 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=15740 $D=0
M1713 767 634 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=20370 $D=0
M1714 164 632 766 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=15740 $D=0
M1715 165 633 767 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=20370 $D=0
M1716 634 766 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=15740 $D=0
M1717 635 767 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=20370 $D=0
M1718 780 533 164 164 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=15380 $D=0
M1719 781 534 165 165 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=20010 $D=0
M1720 636 638 780 164 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=15380 $D=0
M1721 637 639 781 165 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=20010 $D=0
M1722 638 626 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=15740 $D=0
M1723 639 627 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=20370 $D=0
M1724 640 636 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=15740 $D=0
M1725 641 637 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=20370 $D=0
M1726 164 157 640 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=15740 $D=0
M1727 165 634 641 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=20370 $D=0
M1728 643 158 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=15740 $D=0
M1729 644 642 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=20370 $D=0
M1730 642 640 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=15740 $D=0
M1731 159 641 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=20370 $D=0
M1732 164 643 642 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=15740 $D=0
M1733 165 644 159 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=20370 $D=0
M1734 646 645 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=15740 $D=0
M1735 647 160 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=20370 $D=0
M1736 164 650 648 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=15740 $D=0
M1737 165 651 649 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=20370 $D=0
M1738 652 117 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=15740 $D=0
M1739 653 118 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=20370 $D=0
M1740 650 117 645 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=15740 $D=0
M1741 651 118 160 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=20370 $D=0
M1742 646 652 650 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=15740 $D=0
M1743 647 653 651 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=20370 $D=0
M1744 654 648 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=15740 $D=0
M1745 655 649 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=20370 $D=0
M1746 161 648 6 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=15740 $D=0
M1747 645 649 7 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=20370 $D=0
M1748 117 654 161 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=15740 $D=0
M1749 118 655 645 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=20370 $D=0
M1750 656 161 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=15740 $D=0
M1751 657 645 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=20370 $D=0
M1752 658 648 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=15740 $D=0
M1753 659 649 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=20370 $D=0
M1754 195 648 656 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=15740 $D=0
M1755 196 649 657 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=20370 $D=0
M1756 6 658 195 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=15740 $D=0
M1757 7 659 196 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=20370 $D=0
M1758 660 162 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=15740 $D=0
M1759 661 162 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=20370 $D=0
M1760 662 162 195 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=15740 $D=0
M1761 663 162 196 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=20370 $D=0
M1762 14 660 662 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=15740 $D=0
M1763 15 661 663 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=20370 $D=0
M1764 664 163 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=15740 $D=0
M1765 665 163 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=20370 $D=0
M1766 163 163 662 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=15740 $D=0
M1767 163 163 663 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=20370 $D=0
M1768 6 664 163 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=15740 $D=0
M1769 7 665 163 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=20370 $D=0
M1770 666 113 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=15740 $D=0
M1771 667 113 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=20370 $D=0
M1772 164 666 668 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=15740 $D=0
M1773 165 667 669 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=20370 $D=0
M1774 670 113 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=15740 $D=0
M1775 671 113 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=20370 $D=0
M1776 672 668 163 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=15740 $D=0
M1777 673 669 163 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=20370 $D=0
M1778 164 672 768 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=15740 $D=0
M1779 165 673 769 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=20370 $D=0
M1780 674 768 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=15740 $D=0
M1781 675 769 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=20370 $D=0
M1782 672 666 674 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=15740 $D=0
M1783 673 667 675 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=20370 $D=0
M1784 676 670 674 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=15740 $D=0
M1785 677 671 675 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=20370 $D=0
M1786 164 680 678 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=15740 $D=0
M1787 165 681 679 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=20370 $D=0
M1788 680 113 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=15740 $D=0
M1789 681 113 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=20370 $D=0
M1790 770 676 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=15740 $D=0
M1791 771 677 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=20370 $D=0
M1792 682 680 770 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=15740 $D=0
M1793 683 681 771 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=20370 $D=0
M1794 164 682 117 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=15740 $D=0
M1795 165 683 118 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=20370 $D=0
M1796 772 117 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=15740 $D=0
M1797 773 118 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=20370 $D=0
M1798 682 678 772 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=15740 $D=0
M1799 683 679 773 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=20370 $D=0
.ENDS
***************************************
.SUBCKT ICV_41 1 2 3 4 5 6 7 8 9 11 12 13 14 15 16 17 18 19 20 21
+ 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41
+ 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61
+ 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81
+ 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101
+ 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121
+ 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141
+ 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161
+ 162 163 164 165 166 167 168 169 170 171 172 173 174
** N=1124 EP=173 IP=2241 FDC=2700
M0 177 1 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=600 $D=1
M1 178 1 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=5230 $D=1
M2 179 1 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=9860 $D=1
M3 180 177 2 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=600 $D=1
M4 181 178 3 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=5230 $D=1
M5 182 179 4 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=9860 $D=1
M6 7 1 180 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=600 $D=1
M7 8 1 181 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=5230 $D=1
M8 9 1 182 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=9860 $D=1
M9 183 177 5 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=600 $D=1
M10 184 178 5 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=5230 $D=1
M11 185 179 5 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=9860 $D=1
M12 6 1 183 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=600 $D=1
M13 6 1 184 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=5230 $D=1
M14 6 1 185 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=9860 $D=1
M15 186 177 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=600 $D=1
M16 187 178 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=5230 $D=1
M17 188 179 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=9860 $D=1
M18 7 1 186 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=600 $D=1
M19 8 1 187 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=5230 $D=1
M20 9 1 188 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=9860 $D=1
M21 192 189 186 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=600 $D=1
M22 193 190 187 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=5230 $D=1
M23 194 191 188 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=9860 $D=1
M24 189 11 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=600 $D=1
M25 190 11 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=5230 $D=1
M26 191 11 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=9860 $D=1
M27 195 189 183 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=600 $D=1
M28 196 190 184 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=5230 $D=1
M29 197 191 185 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=9860 $D=1
M30 180 11 195 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=600 $D=1
M31 181 11 196 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=5230 $D=1
M32 182 11 197 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=9860 $D=1
M33 198 12 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=600 $D=1
M34 199 12 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=5230 $D=1
M35 200 12 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=9860 $D=1
M36 201 198 195 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=600 $D=1
M37 202 199 196 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=5230 $D=1
M38 203 200 197 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=9860 $D=1
M39 192 12 201 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=600 $D=1
M40 193 12 202 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=5230 $D=1
M41 194 12 203 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=9860 $D=1
M42 204 13 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=600 $D=1
M43 205 13 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=5230 $D=1
M44 206 13 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=9860 $D=1
M45 207 204 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=600 $D=1
M46 208 205 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=5230 $D=1
M47 209 206 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=9860 $D=1
M48 14 13 207 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=600 $D=1
M49 15 13 208 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=5230 $D=1
M50 16 13 209 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=9860 $D=1
M51 210 204 17 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=600 $D=1
M52 211 205 18 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=5230 $D=1
M53 212 206 19 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=9860 $D=1
M54 213 13 210 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=600 $D=1
M55 214 13 211 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=5230 $D=1
M56 215 13 212 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=9860 $D=1
M57 219 204 216 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=600 $D=1
M58 220 205 217 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=5230 $D=1
M59 221 206 218 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=9860 $D=1
M60 201 13 219 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=600 $D=1
M61 202 13 220 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=5230 $D=1
M62 203 13 221 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=9860 $D=1
M63 225 222 219 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=600 $D=1
M64 226 223 220 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=5230 $D=1
M65 227 224 221 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=9860 $D=1
M66 222 20 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=600 $D=1
M67 223 20 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=5230 $D=1
M68 224 20 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=9860 $D=1
M69 228 222 210 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=600 $D=1
M70 229 223 211 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=5230 $D=1
M71 230 224 212 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=9860 $D=1
M72 207 20 228 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=600 $D=1
M73 208 20 229 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=5230 $D=1
M74 209 20 230 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=9860 $D=1
M75 231 21 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=600 $D=1
M76 232 21 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=5230 $D=1
M77 233 21 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=9860 $D=1
M78 234 231 228 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=600 $D=1
M79 235 232 229 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=5230 $D=1
M80 236 233 230 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=9860 $D=1
M81 225 21 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=600 $D=1
M82 226 21 235 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=5230 $D=1
M83 227 21 236 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=9860 $D=1
M84 7 22 237 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=600 $D=1
M85 8 22 238 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=5230 $D=1
M86 9 22 239 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=9860 $D=1
M87 240 23 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=600 $D=1
M88 241 23 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=5230 $D=1
M89 242 23 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=9860 $D=1
M90 243 22 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=600 $D=1
M91 244 22 235 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=5230 $D=1
M92 245 22 236 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=9860 $D=1
M93 7 243 957 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=600 $D=1
M94 8 244 958 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=5230 $D=1
M95 9 245 959 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=9860 $D=1
M96 246 957 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=600 $D=1
M97 247 958 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=5230 $D=1
M98 248 959 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=9860 $D=1
M99 243 237 246 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=600 $D=1
M100 244 238 247 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=5230 $D=1
M101 245 239 248 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=9860 $D=1
M102 246 23 249 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=600 $D=1
M103 247 23 250 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=5230 $D=1
M104 248 23 251 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=9860 $D=1
M105 255 24 246 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=600 $D=1
M106 256 24 247 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=5230 $D=1
M107 257 24 248 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=9860 $D=1
M108 252 24 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=600 $D=1
M109 253 24 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=5230 $D=1
M110 254 24 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=9860 $D=1
M111 7 25 258 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=600 $D=1
M112 8 25 259 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=5230 $D=1
M113 9 25 260 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=9860 $D=1
M114 261 26 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=600 $D=1
M115 262 26 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=5230 $D=1
M116 263 26 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=9860 $D=1
M117 264 25 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=600 $D=1
M118 265 25 235 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=5230 $D=1
M119 266 25 236 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=9860 $D=1
M120 7 264 960 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=600 $D=1
M121 8 265 961 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=5230 $D=1
M122 9 266 962 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=9860 $D=1
M123 267 960 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=600 $D=1
M124 268 961 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=5230 $D=1
M125 269 962 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=9860 $D=1
M126 264 258 267 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=600 $D=1
M127 265 259 268 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=5230 $D=1
M128 266 260 269 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=9860 $D=1
M129 267 26 249 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=600 $D=1
M130 268 26 250 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=5230 $D=1
M131 269 26 251 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=9860 $D=1
M132 255 27 267 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=600 $D=1
M133 256 27 268 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=5230 $D=1
M134 257 27 269 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=9860 $D=1
M135 270 27 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=600 $D=1
M136 271 27 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=5230 $D=1
M137 272 27 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=9860 $D=1
M138 7 28 273 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=600 $D=1
M139 8 28 274 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=5230 $D=1
M140 9 28 275 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=9860 $D=1
M141 276 29 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=600 $D=1
M142 277 29 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=5230 $D=1
M143 278 29 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=9860 $D=1
M144 279 28 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=600 $D=1
M145 280 28 235 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=5230 $D=1
M146 281 28 236 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=9860 $D=1
M147 7 279 963 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=600 $D=1
M148 8 280 964 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=5230 $D=1
M149 9 281 965 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=9860 $D=1
M150 282 963 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=600 $D=1
M151 283 964 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=5230 $D=1
M152 284 965 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=9860 $D=1
M153 279 273 282 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=600 $D=1
M154 280 274 283 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=5230 $D=1
M155 281 275 284 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=9860 $D=1
M156 282 29 249 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=600 $D=1
M157 283 29 250 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=5230 $D=1
M158 284 29 251 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=9860 $D=1
M159 255 30 282 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=600 $D=1
M160 256 30 283 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=5230 $D=1
M161 257 30 284 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=9860 $D=1
M162 285 30 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=600 $D=1
M163 286 30 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=5230 $D=1
M164 287 30 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=9860 $D=1
M165 7 31 288 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=600 $D=1
M166 8 31 289 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=5230 $D=1
M167 9 31 290 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=9860 $D=1
M168 291 32 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=600 $D=1
M169 292 32 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=5230 $D=1
M170 293 32 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=9860 $D=1
M171 294 31 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=600 $D=1
M172 295 31 235 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=5230 $D=1
M173 296 31 236 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=9860 $D=1
M174 7 294 966 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=600 $D=1
M175 8 295 967 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=5230 $D=1
M176 9 296 968 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=9860 $D=1
M177 297 966 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=600 $D=1
M178 298 967 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=5230 $D=1
M179 299 968 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=9860 $D=1
M180 294 288 297 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=600 $D=1
M181 295 289 298 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=5230 $D=1
M182 296 290 299 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=9860 $D=1
M183 297 32 249 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=600 $D=1
M184 298 32 250 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=5230 $D=1
M185 299 32 251 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=9860 $D=1
M186 255 33 297 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=600 $D=1
M187 256 33 298 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=5230 $D=1
M188 257 33 299 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=9860 $D=1
M189 300 33 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=600 $D=1
M190 301 33 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=5230 $D=1
M191 302 33 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=9860 $D=1
M192 7 34 303 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=600 $D=1
M193 8 34 304 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=5230 $D=1
M194 9 34 305 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=9860 $D=1
M195 306 35 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=600 $D=1
M196 307 35 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=5230 $D=1
M197 308 35 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=9860 $D=1
M198 309 34 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=600 $D=1
M199 310 34 235 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=5230 $D=1
M200 311 34 236 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=9860 $D=1
M201 7 309 969 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=600 $D=1
M202 8 310 970 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=5230 $D=1
M203 9 311 971 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=9860 $D=1
M204 312 969 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=600 $D=1
M205 313 970 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=5230 $D=1
M206 314 971 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=9860 $D=1
M207 309 303 312 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=600 $D=1
M208 310 304 313 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=5230 $D=1
M209 311 305 314 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=9860 $D=1
M210 312 35 249 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=600 $D=1
M211 313 35 250 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=5230 $D=1
M212 314 35 251 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=9860 $D=1
M213 255 36 312 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=600 $D=1
M214 256 36 313 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=5230 $D=1
M215 257 36 314 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=9860 $D=1
M216 315 36 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=600 $D=1
M217 316 36 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=5230 $D=1
M218 317 36 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=9860 $D=1
M219 7 37 318 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=600 $D=1
M220 8 37 319 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=5230 $D=1
M221 9 37 320 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=9860 $D=1
M222 321 38 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=600 $D=1
M223 322 38 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=5230 $D=1
M224 323 38 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=9860 $D=1
M225 324 37 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=600 $D=1
M226 325 37 235 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=5230 $D=1
M227 326 37 236 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=9860 $D=1
M228 7 324 972 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=600 $D=1
M229 8 325 973 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=5230 $D=1
M230 9 326 974 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=9860 $D=1
M231 327 972 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=600 $D=1
M232 328 973 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=5230 $D=1
M233 329 974 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=9860 $D=1
M234 324 318 327 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=600 $D=1
M235 325 319 328 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=5230 $D=1
M236 326 320 329 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=9860 $D=1
M237 327 38 249 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=600 $D=1
M238 328 38 250 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=5230 $D=1
M239 329 38 251 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=9860 $D=1
M240 255 39 327 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=600 $D=1
M241 256 39 328 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=5230 $D=1
M242 257 39 329 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=9860 $D=1
M243 330 39 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=600 $D=1
M244 331 39 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=5230 $D=1
M245 332 39 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=9860 $D=1
M246 7 40 333 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=600 $D=1
M247 8 40 334 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=5230 $D=1
M248 9 40 335 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=9860 $D=1
M249 336 41 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=600 $D=1
M250 337 41 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=5230 $D=1
M251 338 41 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=9860 $D=1
M252 339 40 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=600 $D=1
M253 340 40 235 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=5230 $D=1
M254 341 40 236 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=9860 $D=1
M255 7 339 975 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=600 $D=1
M256 8 340 976 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=5230 $D=1
M257 9 341 977 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=9860 $D=1
M258 342 975 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=600 $D=1
M259 343 976 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=5230 $D=1
M260 344 977 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=9860 $D=1
M261 339 333 342 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=600 $D=1
M262 340 334 343 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=5230 $D=1
M263 341 335 344 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=9860 $D=1
M264 342 41 249 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=600 $D=1
M265 343 41 250 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=5230 $D=1
M266 344 41 251 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=9860 $D=1
M267 255 42 342 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=600 $D=1
M268 256 42 343 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=5230 $D=1
M269 257 42 344 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=9860 $D=1
M270 345 42 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=600 $D=1
M271 346 42 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=5230 $D=1
M272 347 42 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=9860 $D=1
M273 7 43 348 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=600 $D=1
M274 8 43 349 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=5230 $D=1
M275 9 43 350 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=9860 $D=1
M276 351 44 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=600 $D=1
M277 352 44 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=5230 $D=1
M278 353 44 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=9860 $D=1
M279 354 43 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=600 $D=1
M280 355 43 235 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=5230 $D=1
M281 356 43 236 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=9860 $D=1
M282 7 354 978 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=600 $D=1
M283 8 355 979 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=5230 $D=1
M284 9 356 980 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=9860 $D=1
M285 357 978 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=600 $D=1
M286 358 979 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=5230 $D=1
M287 359 980 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=9860 $D=1
M288 354 348 357 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=600 $D=1
M289 355 349 358 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=5230 $D=1
M290 356 350 359 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=9860 $D=1
M291 357 44 249 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=600 $D=1
M292 358 44 250 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=5230 $D=1
M293 359 44 251 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=9860 $D=1
M294 255 45 357 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=600 $D=1
M295 256 45 358 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=5230 $D=1
M296 257 45 359 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=9860 $D=1
M297 360 45 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=600 $D=1
M298 361 45 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=5230 $D=1
M299 362 45 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=9860 $D=1
M300 7 46 363 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=600 $D=1
M301 8 46 364 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=5230 $D=1
M302 9 46 365 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=9860 $D=1
M303 366 47 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=600 $D=1
M304 367 47 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=5230 $D=1
M305 368 47 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=9860 $D=1
M306 369 46 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=600 $D=1
M307 370 46 235 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=5230 $D=1
M308 371 46 236 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=9860 $D=1
M309 7 369 981 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=600 $D=1
M310 8 370 982 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=5230 $D=1
M311 9 371 983 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=9860 $D=1
M312 372 981 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=600 $D=1
M313 373 982 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=5230 $D=1
M314 374 983 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=9860 $D=1
M315 369 363 372 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=600 $D=1
M316 370 364 373 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=5230 $D=1
M317 371 365 374 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=9860 $D=1
M318 372 47 249 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=600 $D=1
M319 373 47 250 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=5230 $D=1
M320 374 47 251 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=9860 $D=1
M321 255 48 372 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=600 $D=1
M322 256 48 373 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=5230 $D=1
M323 257 48 374 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=9860 $D=1
M324 375 48 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=600 $D=1
M325 376 48 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=5230 $D=1
M326 377 48 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=9860 $D=1
M327 7 49 378 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=600 $D=1
M328 8 49 379 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=5230 $D=1
M329 9 49 380 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=9860 $D=1
M330 381 50 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=600 $D=1
M331 382 50 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=5230 $D=1
M332 383 50 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=9860 $D=1
M333 384 49 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=600 $D=1
M334 385 49 235 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=5230 $D=1
M335 386 49 236 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=9860 $D=1
M336 7 384 984 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=600 $D=1
M337 8 385 985 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=5230 $D=1
M338 9 386 986 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=9860 $D=1
M339 387 984 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=600 $D=1
M340 388 985 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=5230 $D=1
M341 389 986 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=9860 $D=1
M342 384 378 387 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=600 $D=1
M343 385 379 388 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=5230 $D=1
M344 386 380 389 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=9860 $D=1
M345 387 50 249 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=600 $D=1
M346 388 50 250 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=5230 $D=1
M347 389 50 251 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=9860 $D=1
M348 255 51 387 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=600 $D=1
M349 256 51 388 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=5230 $D=1
M350 257 51 389 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=9860 $D=1
M351 390 51 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=600 $D=1
M352 391 51 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=5230 $D=1
M353 392 51 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=9860 $D=1
M354 7 52 393 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=600 $D=1
M355 8 52 394 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=5230 $D=1
M356 9 52 395 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=9860 $D=1
M357 396 53 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=600 $D=1
M358 397 53 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=5230 $D=1
M359 398 53 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=9860 $D=1
M360 399 52 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=600 $D=1
M361 400 52 235 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=5230 $D=1
M362 401 52 236 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=9860 $D=1
M363 7 399 987 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=600 $D=1
M364 8 400 988 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=5230 $D=1
M365 9 401 989 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=9860 $D=1
M366 402 987 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=600 $D=1
M367 403 988 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=5230 $D=1
M368 404 989 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=9860 $D=1
M369 399 393 402 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=600 $D=1
M370 400 394 403 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=5230 $D=1
M371 401 395 404 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=9860 $D=1
M372 402 53 249 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=600 $D=1
M373 403 53 250 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=5230 $D=1
M374 404 53 251 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=9860 $D=1
M375 255 54 402 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=600 $D=1
M376 256 54 403 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=5230 $D=1
M377 257 54 404 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=9860 $D=1
M378 405 54 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=600 $D=1
M379 406 54 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=5230 $D=1
M380 407 54 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=9860 $D=1
M381 7 55 408 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=600 $D=1
M382 8 55 409 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=5230 $D=1
M383 9 55 410 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=9860 $D=1
M384 411 56 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=600 $D=1
M385 412 56 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=5230 $D=1
M386 413 56 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=9860 $D=1
M387 414 55 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=600 $D=1
M388 415 55 235 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=5230 $D=1
M389 416 55 236 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=9860 $D=1
M390 7 414 990 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=600 $D=1
M391 8 415 991 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=5230 $D=1
M392 9 416 992 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=9860 $D=1
M393 417 990 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=600 $D=1
M394 418 991 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=5230 $D=1
M395 419 992 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=9860 $D=1
M396 414 408 417 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=600 $D=1
M397 415 409 418 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=5230 $D=1
M398 416 410 419 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=9860 $D=1
M399 417 56 249 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=600 $D=1
M400 418 56 250 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=5230 $D=1
M401 419 56 251 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=9860 $D=1
M402 255 57 417 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=600 $D=1
M403 256 57 418 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=5230 $D=1
M404 257 57 419 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=9860 $D=1
M405 420 57 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=600 $D=1
M406 421 57 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=5230 $D=1
M407 422 57 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=9860 $D=1
M408 7 58 423 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=600 $D=1
M409 8 58 424 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=5230 $D=1
M410 9 58 425 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=9860 $D=1
M411 426 59 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=600 $D=1
M412 427 59 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=5230 $D=1
M413 428 59 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=9860 $D=1
M414 429 58 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=600 $D=1
M415 430 58 235 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=5230 $D=1
M416 431 58 236 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=9860 $D=1
M417 7 429 993 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=600 $D=1
M418 8 430 994 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=5230 $D=1
M419 9 431 995 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=9860 $D=1
M420 432 993 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=600 $D=1
M421 433 994 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=5230 $D=1
M422 434 995 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=9860 $D=1
M423 429 423 432 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=600 $D=1
M424 430 424 433 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=5230 $D=1
M425 431 425 434 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=9860 $D=1
M426 432 59 249 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=600 $D=1
M427 433 59 250 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=5230 $D=1
M428 434 59 251 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=9860 $D=1
M429 255 60 432 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=600 $D=1
M430 256 60 433 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=5230 $D=1
M431 257 60 434 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=9860 $D=1
M432 435 60 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=600 $D=1
M433 436 60 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=5230 $D=1
M434 437 60 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=9860 $D=1
M435 7 61 438 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=600 $D=1
M436 8 61 439 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=5230 $D=1
M437 9 61 440 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=9860 $D=1
M438 441 62 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=600 $D=1
M439 442 62 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=5230 $D=1
M440 443 62 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=9860 $D=1
M441 444 61 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=600 $D=1
M442 445 61 235 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=5230 $D=1
M443 446 61 236 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=9860 $D=1
M444 7 444 996 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=600 $D=1
M445 8 445 997 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=5230 $D=1
M446 9 446 998 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=9860 $D=1
M447 447 996 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=600 $D=1
M448 448 997 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=5230 $D=1
M449 449 998 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=9860 $D=1
M450 444 438 447 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=600 $D=1
M451 445 439 448 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=5230 $D=1
M452 446 440 449 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=9860 $D=1
M453 447 62 249 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=600 $D=1
M454 448 62 250 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=5230 $D=1
M455 449 62 251 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=9860 $D=1
M456 255 63 447 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=600 $D=1
M457 256 63 448 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=5230 $D=1
M458 257 63 449 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=9860 $D=1
M459 450 63 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=600 $D=1
M460 451 63 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=5230 $D=1
M461 452 63 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=9860 $D=1
M462 7 64 453 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=600 $D=1
M463 8 64 454 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=5230 $D=1
M464 9 64 455 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=9860 $D=1
M465 456 65 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=600 $D=1
M466 457 65 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=5230 $D=1
M467 458 65 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=9860 $D=1
M468 459 64 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=600 $D=1
M469 460 64 235 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=5230 $D=1
M470 461 64 236 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=9860 $D=1
M471 7 459 999 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=600 $D=1
M472 8 460 1000 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=5230 $D=1
M473 9 461 1001 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=9860 $D=1
M474 462 999 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=600 $D=1
M475 463 1000 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=5230 $D=1
M476 464 1001 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=9860 $D=1
M477 459 453 462 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=600 $D=1
M478 460 454 463 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=5230 $D=1
M479 461 455 464 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=9860 $D=1
M480 462 65 249 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=600 $D=1
M481 463 65 250 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=5230 $D=1
M482 464 65 251 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=9860 $D=1
M483 255 66 462 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=600 $D=1
M484 256 66 463 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=5230 $D=1
M485 257 66 464 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=9860 $D=1
M486 465 66 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=600 $D=1
M487 466 66 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=5230 $D=1
M488 467 66 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=9860 $D=1
M489 7 67 468 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=600 $D=1
M490 8 67 469 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=5230 $D=1
M491 9 67 470 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=9860 $D=1
M492 471 68 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=600 $D=1
M493 472 68 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=5230 $D=1
M494 473 68 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=9860 $D=1
M495 474 67 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=600 $D=1
M496 475 67 235 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=5230 $D=1
M497 476 67 236 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=9860 $D=1
M498 7 474 1002 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=600 $D=1
M499 8 475 1003 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=5230 $D=1
M500 9 476 1004 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=9860 $D=1
M501 477 1002 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=600 $D=1
M502 478 1003 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=5230 $D=1
M503 479 1004 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=9860 $D=1
M504 474 468 477 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=600 $D=1
M505 475 469 478 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=5230 $D=1
M506 476 470 479 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=9860 $D=1
M507 477 68 249 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=600 $D=1
M508 478 68 250 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=5230 $D=1
M509 479 68 251 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=9860 $D=1
M510 255 69 477 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=600 $D=1
M511 256 69 478 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=5230 $D=1
M512 257 69 479 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=9860 $D=1
M513 480 69 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=600 $D=1
M514 481 69 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=5230 $D=1
M515 482 69 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=9860 $D=1
M516 7 70 483 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=600 $D=1
M517 8 70 484 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=5230 $D=1
M518 9 70 485 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=9860 $D=1
M519 486 71 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=600 $D=1
M520 487 71 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=5230 $D=1
M521 488 71 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=9860 $D=1
M522 489 70 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=600 $D=1
M523 490 70 235 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=5230 $D=1
M524 491 70 236 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=9860 $D=1
M525 7 489 1005 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=600 $D=1
M526 8 490 1006 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=5230 $D=1
M527 9 491 1007 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=9860 $D=1
M528 492 1005 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=600 $D=1
M529 493 1006 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=5230 $D=1
M530 494 1007 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=9860 $D=1
M531 489 483 492 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=600 $D=1
M532 490 484 493 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=5230 $D=1
M533 491 485 494 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=9860 $D=1
M534 492 71 249 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=600 $D=1
M535 493 71 250 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=5230 $D=1
M536 494 71 251 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=9860 $D=1
M537 255 72 492 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=600 $D=1
M538 256 72 493 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=5230 $D=1
M539 257 72 494 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=9860 $D=1
M540 495 72 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=600 $D=1
M541 496 72 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=5230 $D=1
M542 497 72 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=9860 $D=1
M543 7 73 498 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=600 $D=1
M544 8 73 499 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=5230 $D=1
M545 9 73 500 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=9860 $D=1
M546 501 74 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=600 $D=1
M547 502 74 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=5230 $D=1
M548 503 74 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=9860 $D=1
M549 504 73 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=600 $D=1
M550 505 73 235 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=5230 $D=1
M551 506 73 236 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=9860 $D=1
M552 7 504 1008 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=600 $D=1
M553 8 505 1009 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=5230 $D=1
M554 9 506 1010 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=9860 $D=1
M555 507 1008 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=600 $D=1
M556 508 1009 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=5230 $D=1
M557 509 1010 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=9860 $D=1
M558 504 498 507 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=600 $D=1
M559 505 499 508 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=5230 $D=1
M560 506 500 509 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=9860 $D=1
M561 507 74 249 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=600 $D=1
M562 508 74 250 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=5230 $D=1
M563 509 74 251 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=9860 $D=1
M564 255 75 507 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=600 $D=1
M565 256 75 508 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=5230 $D=1
M566 257 75 509 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=9860 $D=1
M567 510 75 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=600 $D=1
M568 511 75 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=5230 $D=1
M569 512 75 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=9860 $D=1
M570 7 76 513 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=600 $D=1
M571 8 76 514 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=5230 $D=1
M572 9 76 515 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=9860 $D=1
M573 516 77 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=600 $D=1
M574 517 77 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=5230 $D=1
M575 518 77 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=9860 $D=1
M576 519 76 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=600 $D=1
M577 520 76 235 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=5230 $D=1
M578 521 76 236 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=9860 $D=1
M579 7 519 1011 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=600 $D=1
M580 8 520 1012 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=5230 $D=1
M581 9 521 1013 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=9860 $D=1
M582 522 1011 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=600 $D=1
M583 523 1012 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=5230 $D=1
M584 524 1013 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=9860 $D=1
M585 519 513 522 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=600 $D=1
M586 520 514 523 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=5230 $D=1
M587 521 515 524 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=9860 $D=1
M588 522 77 249 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=600 $D=1
M589 523 77 250 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=5230 $D=1
M590 524 77 251 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=9860 $D=1
M591 255 78 522 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=600 $D=1
M592 256 78 523 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=5230 $D=1
M593 257 78 524 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=9860 $D=1
M594 525 78 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=600 $D=1
M595 526 78 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=5230 $D=1
M596 527 78 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=9860 $D=1
M597 7 79 528 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=600 $D=1
M598 8 79 529 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=5230 $D=1
M599 9 79 530 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=9860 $D=1
M600 531 80 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=600 $D=1
M601 532 80 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=5230 $D=1
M602 533 80 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=9860 $D=1
M603 534 79 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=600 $D=1
M604 535 79 235 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=5230 $D=1
M605 536 79 236 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=9860 $D=1
M606 7 534 1014 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=600 $D=1
M607 8 535 1015 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=5230 $D=1
M608 9 536 1016 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=9860 $D=1
M609 537 1014 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=600 $D=1
M610 538 1015 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=5230 $D=1
M611 539 1016 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=9860 $D=1
M612 534 528 537 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=600 $D=1
M613 535 529 538 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=5230 $D=1
M614 536 530 539 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=9860 $D=1
M615 537 80 249 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=600 $D=1
M616 538 80 250 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=5230 $D=1
M617 539 80 251 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=9860 $D=1
M618 255 81 537 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=600 $D=1
M619 256 81 538 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=5230 $D=1
M620 257 81 539 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=9860 $D=1
M621 540 81 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=600 $D=1
M622 541 81 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=5230 $D=1
M623 542 81 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=9860 $D=1
M624 7 82 543 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=600 $D=1
M625 8 82 544 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=5230 $D=1
M626 9 82 545 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=9860 $D=1
M627 546 83 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=600 $D=1
M628 547 83 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=5230 $D=1
M629 548 83 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=9860 $D=1
M630 549 82 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=600 $D=1
M631 550 82 235 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=5230 $D=1
M632 551 82 236 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=9860 $D=1
M633 7 549 1017 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=600 $D=1
M634 8 550 1018 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=5230 $D=1
M635 9 551 1019 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=9860 $D=1
M636 552 1017 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=600 $D=1
M637 553 1018 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=5230 $D=1
M638 554 1019 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=9860 $D=1
M639 549 543 552 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=600 $D=1
M640 550 544 553 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=5230 $D=1
M641 551 545 554 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=9860 $D=1
M642 552 83 249 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=600 $D=1
M643 553 83 250 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=5230 $D=1
M644 554 83 251 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=9860 $D=1
M645 255 84 552 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=600 $D=1
M646 256 84 553 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=5230 $D=1
M647 257 84 554 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=9860 $D=1
M648 555 84 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=600 $D=1
M649 556 84 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=5230 $D=1
M650 557 84 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=9860 $D=1
M651 7 85 558 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=600 $D=1
M652 8 85 559 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=5230 $D=1
M653 9 85 560 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=9860 $D=1
M654 561 86 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=600 $D=1
M655 562 86 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=5230 $D=1
M656 563 86 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=9860 $D=1
M657 564 85 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=600 $D=1
M658 565 85 235 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=5230 $D=1
M659 566 85 236 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=9860 $D=1
M660 7 564 1020 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=600 $D=1
M661 8 565 1021 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=5230 $D=1
M662 9 566 1022 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=9860 $D=1
M663 567 1020 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=600 $D=1
M664 568 1021 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=5230 $D=1
M665 569 1022 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=9860 $D=1
M666 564 558 567 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=600 $D=1
M667 565 559 568 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=5230 $D=1
M668 566 560 569 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=9860 $D=1
M669 567 86 249 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=600 $D=1
M670 568 86 250 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=5230 $D=1
M671 569 86 251 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=9860 $D=1
M672 255 87 567 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=600 $D=1
M673 256 87 568 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=5230 $D=1
M674 257 87 569 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=9860 $D=1
M675 570 87 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=600 $D=1
M676 571 87 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=5230 $D=1
M677 572 87 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=9860 $D=1
M678 7 88 573 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=600 $D=1
M679 8 88 574 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=5230 $D=1
M680 9 88 575 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=9860 $D=1
M681 576 89 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=600 $D=1
M682 577 89 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=5230 $D=1
M683 578 89 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=9860 $D=1
M684 579 88 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=600 $D=1
M685 580 88 235 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=5230 $D=1
M686 581 88 236 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=9860 $D=1
M687 7 579 1023 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=600 $D=1
M688 8 580 1024 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=5230 $D=1
M689 9 581 1025 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=9860 $D=1
M690 582 1023 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=600 $D=1
M691 583 1024 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=5230 $D=1
M692 584 1025 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=9860 $D=1
M693 579 573 582 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=600 $D=1
M694 580 574 583 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=5230 $D=1
M695 581 575 584 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=9860 $D=1
M696 582 89 249 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=600 $D=1
M697 583 89 250 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=5230 $D=1
M698 584 89 251 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=9860 $D=1
M699 255 90 582 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=600 $D=1
M700 256 90 583 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=5230 $D=1
M701 257 90 584 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=9860 $D=1
M702 585 90 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=600 $D=1
M703 586 90 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=5230 $D=1
M704 587 90 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=9860 $D=1
M705 7 91 588 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=600 $D=1
M706 8 91 589 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=5230 $D=1
M707 9 91 590 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=9860 $D=1
M708 591 92 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=600 $D=1
M709 592 92 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=5230 $D=1
M710 593 92 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=9860 $D=1
M711 594 91 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=600 $D=1
M712 595 91 235 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=5230 $D=1
M713 596 91 236 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=9860 $D=1
M714 7 594 1026 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=600 $D=1
M715 8 595 1027 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=5230 $D=1
M716 9 596 1028 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=9860 $D=1
M717 597 1026 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=600 $D=1
M718 598 1027 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=5230 $D=1
M719 599 1028 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=9860 $D=1
M720 594 588 597 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=600 $D=1
M721 595 589 598 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=5230 $D=1
M722 596 590 599 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=9860 $D=1
M723 597 92 249 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=600 $D=1
M724 598 92 250 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=5230 $D=1
M725 599 92 251 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=9860 $D=1
M726 255 93 597 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=600 $D=1
M727 256 93 598 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=5230 $D=1
M728 257 93 599 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=9860 $D=1
M729 600 93 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=600 $D=1
M730 601 93 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=5230 $D=1
M731 602 93 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=9860 $D=1
M732 7 94 603 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=600 $D=1
M733 8 94 604 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=5230 $D=1
M734 9 94 605 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=9860 $D=1
M735 606 95 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=600 $D=1
M736 607 95 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=5230 $D=1
M737 608 95 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=9860 $D=1
M738 609 94 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=600 $D=1
M739 610 94 235 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=5230 $D=1
M740 611 94 236 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=9860 $D=1
M741 7 609 1029 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=600 $D=1
M742 8 610 1030 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=5230 $D=1
M743 9 611 1031 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=9860 $D=1
M744 612 1029 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=600 $D=1
M745 613 1030 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=5230 $D=1
M746 614 1031 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=9860 $D=1
M747 609 603 612 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=600 $D=1
M748 610 604 613 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=5230 $D=1
M749 611 605 614 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=9860 $D=1
M750 612 95 249 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=600 $D=1
M751 613 95 250 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=5230 $D=1
M752 614 95 251 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=9860 $D=1
M753 255 96 612 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=600 $D=1
M754 256 96 613 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=5230 $D=1
M755 257 96 614 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=9860 $D=1
M756 615 96 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=600 $D=1
M757 616 96 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=5230 $D=1
M758 617 96 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=9860 $D=1
M759 7 97 618 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=600 $D=1
M760 8 97 619 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=5230 $D=1
M761 9 97 620 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=9860 $D=1
M762 621 98 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=600 $D=1
M763 622 98 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=5230 $D=1
M764 623 98 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=9860 $D=1
M765 624 97 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=600 $D=1
M766 625 97 235 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=5230 $D=1
M767 626 97 236 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=9860 $D=1
M768 7 624 1032 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=600 $D=1
M769 8 625 1033 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=5230 $D=1
M770 9 626 1034 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=9860 $D=1
M771 627 1032 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=600 $D=1
M772 628 1033 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=5230 $D=1
M773 629 1034 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=9860 $D=1
M774 624 618 627 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=600 $D=1
M775 625 619 628 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=5230 $D=1
M776 626 620 629 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=9860 $D=1
M777 627 98 249 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=600 $D=1
M778 628 98 250 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=5230 $D=1
M779 629 98 251 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=9860 $D=1
M780 255 99 627 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=600 $D=1
M781 256 99 628 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=5230 $D=1
M782 257 99 629 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=9860 $D=1
M783 630 99 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=600 $D=1
M784 631 99 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=5230 $D=1
M785 632 99 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=9860 $D=1
M786 7 100 633 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=600 $D=1
M787 8 100 634 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=5230 $D=1
M788 9 100 635 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=9860 $D=1
M789 636 101 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=600 $D=1
M790 637 101 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=5230 $D=1
M791 638 101 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=9860 $D=1
M792 639 100 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=600 $D=1
M793 640 100 235 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=5230 $D=1
M794 641 100 236 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=9860 $D=1
M795 7 639 1035 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=600 $D=1
M796 8 640 1036 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=5230 $D=1
M797 9 641 1037 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=9860 $D=1
M798 642 1035 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=600 $D=1
M799 643 1036 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=5230 $D=1
M800 644 1037 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=9860 $D=1
M801 639 633 642 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=600 $D=1
M802 640 634 643 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=5230 $D=1
M803 641 635 644 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=9860 $D=1
M804 642 101 249 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=600 $D=1
M805 643 101 250 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=5230 $D=1
M806 644 101 251 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=9860 $D=1
M807 255 102 642 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=600 $D=1
M808 256 102 643 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=5230 $D=1
M809 257 102 644 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=9860 $D=1
M810 645 102 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=600 $D=1
M811 646 102 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=5230 $D=1
M812 647 102 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=9860 $D=1
M813 7 103 648 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=600 $D=1
M814 8 103 649 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=5230 $D=1
M815 9 103 650 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=9860 $D=1
M816 651 104 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=600 $D=1
M817 652 104 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=5230 $D=1
M818 653 104 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=9860 $D=1
M819 654 103 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=600 $D=1
M820 655 103 235 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=5230 $D=1
M821 656 103 236 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=9860 $D=1
M822 7 654 1038 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=600 $D=1
M823 8 655 1039 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=5230 $D=1
M824 9 656 1040 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=9860 $D=1
M825 657 1038 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=600 $D=1
M826 658 1039 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=5230 $D=1
M827 659 1040 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=9860 $D=1
M828 654 648 657 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=600 $D=1
M829 655 649 658 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=5230 $D=1
M830 656 650 659 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=9860 $D=1
M831 657 104 249 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=600 $D=1
M832 658 104 250 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=5230 $D=1
M833 659 104 251 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=9860 $D=1
M834 255 105 657 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=600 $D=1
M835 256 105 658 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=5230 $D=1
M836 257 105 659 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=9860 $D=1
M837 660 105 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=600 $D=1
M838 661 105 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=5230 $D=1
M839 662 105 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=9860 $D=1
M840 7 106 663 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=600 $D=1
M841 8 106 664 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=5230 $D=1
M842 9 106 665 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=9860 $D=1
M843 666 107 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=600 $D=1
M844 667 107 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=5230 $D=1
M845 668 107 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=9860 $D=1
M846 669 106 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=600 $D=1
M847 670 106 235 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=5230 $D=1
M848 671 106 236 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=9860 $D=1
M849 7 669 1041 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=600 $D=1
M850 8 670 1042 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=5230 $D=1
M851 9 671 1043 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=9860 $D=1
M852 672 1041 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=600 $D=1
M853 673 1042 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=5230 $D=1
M854 674 1043 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=9860 $D=1
M855 669 663 672 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=600 $D=1
M856 670 664 673 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=5230 $D=1
M857 671 665 674 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=9860 $D=1
M858 672 107 249 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=600 $D=1
M859 673 107 250 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=5230 $D=1
M860 674 107 251 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=9860 $D=1
M861 255 108 672 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=600 $D=1
M862 256 108 673 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=5230 $D=1
M863 257 108 674 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=9860 $D=1
M864 675 108 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=600 $D=1
M865 676 108 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=5230 $D=1
M866 677 108 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=9860 $D=1
M867 7 109 678 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=600 $D=1
M868 8 109 679 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=5230 $D=1
M869 9 109 680 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=9860 $D=1
M870 681 110 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=600 $D=1
M871 682 110 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=5230 $D=1
M872 683 110 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=9860 $D=1
M873 684 109 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=600 $D=1
M874 685 109 235 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=5230 $D=1
M875 686 109 236 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=9860 $D=1
M876 7 684 1044 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=600 $D=1
M877 8 685 1045 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=5230 $D=1
M878 9 686 1046 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=9860 $D=1
M879 687 1044 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=600 $D=1
M880 688 1045 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=5230 $D=1
M881 689 1046 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=9860 $D=1
M882 684 678 687 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=600 $D=1
M883 685 679 688 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=5230 $D=1
M884 686 680 689 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=9860 $D=1
M885 687 110 249 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=600 $D=1
M886 688 110 250 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=5230 $D=1
M887 689 110 251 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=9860 $D=1
M888 255 111 687 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=600 $D=1
M889 256 111 688 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=5230 $D=1
M890 257 111 689 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=9860 $D=1
M891 690 111 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=600 $D=1
M892 691 111 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=5230 $D=1
M893 692 111 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=9860 $D=1
M894 7 112 693 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=600 $D=1
M895 8 112 694 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=5230 $D=1
M896 9 112 695 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=9860 $D=1
M897 696 113 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=600 $D=1
M898 697 113 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=5230 $D=1
M899 698 113 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=9860 $D=1
M900 699 112 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=600 $D=1
M901 700 112 235 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=5230 $D=1
M902 701 112 236 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=9860 $D=1
M903 7 699 1047 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=600 $D=1
M904 8 700 1048 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=5230 $D=1
M905 9 701 1049 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=9860 $D=1
M906 702 1047 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=600 $D=1
M907 703 1048 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=5230 $D=1
M908 704 1049 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=9860 $D=1
M909 699 693 702 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=600 $D=1
M910 700 694 703 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=5230 $D=1
M911 701 695 704 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=9860 $D=1
M912 702 113 249 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=600 $D=1
M913 703 113 250 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=5230 $D=1
M914 704 113 251 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=9860 $D=1
M915 255 114 702 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=600 $D=1
M916 256 114 703 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=5230 $D=1
M917 257 114 704 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=9860 $D=1
M918 705 114 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=600 $D=1
M919 706 114 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=5230 $D=1
M920 707 114 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=9860 $D=1
M921 7 115 708 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=600 $D=1
M922 8 115 709 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=5230 $D=1
M923 9 115 710 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=9860 $D=1
M924 711 116 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=600 $D=1
M925 712 116 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=5230 $D=1
M926 713 116 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=9860 $D=1
M927 7 116 249 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=600 $D=1
M928 8 116 250 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=5230 $D=1
M929 9 116 251 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=9860 $D=1
M930 255 115 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=600 $D=1
M931 256 115 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=5230 $D=1
M932 257 115 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=9860 $D=1
M933 7 717 714 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=600 $D=1
M934 8 718 715 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=5230 $D=1
M935 9 719 716 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=9860 $D=1
M936 717 117 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=600 $D=1
M937 718 117 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=5230 $D=1
M938 719 117 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=9860 $D=1
M939 1050 249 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=600 $D=1
M940 1051 250 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=5230 $D=1
M941 1052 251 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=9860 $D=1
M942 720 714 1050 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=600 $D=1
M943 721 715 1051 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=5230 $D=1
M944 722 716 1052 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=9860 $D=1
M945 7 720 118 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=600 $D=1
M946 8 721 723 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=5230 $D=1
M947 9 722 724 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=9860 $D=1
M948 1053 118 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=600 $D=1
M949 1054 723 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=5230 $D=1
M950 1055 724 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=9860 $D=1
M951 720 717 1053 7 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=600 $D=1
M952 721 718 1054 8 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=5230 $D=1
M953 722 719 1055 9 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=9860 $D=1
M954 7 728 725 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=600 $D=1
M955 8 729 726 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=5230 $D=1
M956 9 730 727 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=9860 $D=1
M957 728 117 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=600 $D=1
M958 729 117 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=5230 $D=1
M959 730 117 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=9860 $D=1
M960 1056 255 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=600 $D=1
M961 1057 256 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=5230 $D=1
M962 1058 257 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=9860 $D=1
M963 731 725 1056 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=600 $D=1
M964 732 726 1057 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=5230 $D=1
M965 733 727 1058 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=9860 $D=1
M966 7 731 119 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=600 $D=1
M967 8 732 120 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=5230 $D=1
M968 9 733 121 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=9860 $D=1
M969 1059 119 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=600 $D=1
M970 1060 120 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=5230 $D=1
M971 1061 121 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=9860 $D=1
M972 731 728 1059 7 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=600 $D=1
M973 732 729 1060 8 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=5230 $D=1
M974 733 730 1061 9 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=9860 $D=1
M975 734 122 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=600 $D=1
M976 735 122 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=5230 $D=1
M977 736 122 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=9860 $D=1
M978 737 734 118 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=600 $D=1
M979 738 735 723 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=5230 $D=1
M980 739 736 724 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=9860 $D=1
M981 123 122 737 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=600 $D=1
M982 124 122 738 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=5230 $D=1
M983 125 122 739 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=9860 $D=1
M984 740 126 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=600 $D=1
M985 741 126 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=5230 $D=1
M986 742 126 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=9860 $D=1
M987 743 740 119 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=600 $D=1
M988 744 741 120 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=5230 $D=1
M989 745 742 121 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=9860 $D=1
M990 1062 126 743 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=600 $D=1
M991 1063 126 744 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=5230 $D=1
M992 1064 126 745 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=9860 $D=1
M993 7 119 1062 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=600 $D=1
M994 8 120 1063 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=5230 $D=1
M995 9 121 1064 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=9860 $D=1
M996 746 127 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=600 $D=1
M997 747 127 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=5230 $D=1
M998 748 127 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=9860 $D=1
M999 749 746 743 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=600 $D=1
M1000 750 747 744 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=5230 $D=1
M1001 751 748 745 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=9860 $D=1
M1002 14 127 749 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=600 $D=1
M1003 15 127 750 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=5230 $D=1
M1004 16 127 751 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=9860 $D=1
M1005 755 752 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=600 $D=1
M1006 756 753 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=5230 $D=1
M1007 757 754 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=9860 $D=1
M1008 7 761 758 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=600 $D=1
M1009 8 762 759 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=5230 $D=1
M1010 9 763 760 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=9860 $D=1
M1011 764 737 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=600 $D=1
M1012 765 738 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=5230 $D=1
M1013 766 739 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=9860 $D=1
M1014 761 764 752 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=600 $D=1
M1015 762 765 753 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=5230 $D=1
M1016 763 766 754 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=9860 $D=1
M1017 755 737 761 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=600 $D=1
M1018 756 738 762 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=5230 $D=1
M1019 757 739 763 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=9860 $D=1
M1020 767 758 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=600 $D=1
M1021 768 759 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=5230 $D=1
M1022 769 760 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=9860 $D=1
M1023 770 767 749 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=600 $D=1
M1024 771 768 750 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=5230 $D=1
M1025 772 769 751 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=9860 $D=1
M1026 737 758 770 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=600 $D=1
M1027 738 759 771 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=5230 $D=1
M1028 739 760 772 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=9860 $D=1
M1029 773 770 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=600 $D=1
M1030 774 771 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=5230 $D=1
M1031 775 772 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=9860 $D=1
M1032 776 758 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=600 $D=1
M1033 777 759 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=5230 $D=1
M1034 778 760 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=9860 $D=1
M1035 779 776 773 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=600 $D=1
M1036 780 777 774 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=5230 $D=1
M1037 781 778 775 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=9860 $D=1
M1038 749 758 779 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=600 $D=1
M1039 750 759 780 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=5230 $D=1
M1040 751 760 781 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=9860 $D=1
M1041 782 737 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=600 $D=1
M1042 783 738 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=5230 $D=1
M1043 784 739 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=9860 $D=1
M1044 7 749 782 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=600 $D=1
M1045 8 750 783 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=5230 $D=1
M1046 9 751 784 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=9860 $D=1
M1047 785 779 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=600 $D=1
M1048 786 780 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=5230 $D=1
M1049 787 781 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=9860 $D=1
M1050 1107 737 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=600 $D=1
M1051 1108 738 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=5230 $D=1
M1052 1109 739 9 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=9860 $D=1
M1053 788 749 1107 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=600 $D=1
M1054 789 750 1108 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=5230 $D=1
M1055 790 751 1109 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=9860 $D=1
M1056 1110 737 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=600 $D=1
M1057 1111 738 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=5230 $D=1
M1058 1112 739 9 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=9860 $D=1
M1059 791 749 1110 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=600 $D=1
M1060 792 750 1111 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=5230 $D=1
M1061 793 751 1112 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=9860 $D=1
M1062 797 737 794 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=600 $D=1
M1063 798 738 795 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=5230 $D=1
M1064 799 739 796 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=9860 $D=1
M1065 794 749 797 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=600 $D=1
M1066 795 750 798 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=5230 $D=1
M1067 796 751 799 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=9860 $D=1
M1068 7 791 794 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=600 $D=1
M1069 8 792 795 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=5230 $D=1
M1070 9 793 796 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=9860 $D=1
M1071 800 131 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=600 $D=1
M1072 801 131 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=5230 $D=1
M1073 802 131 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=9860 $D=1
M1074 803 800 782 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=600 $D=1
M1075 804 801 783 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=5230 $D=1
M1076 805 802 784 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=9860 $D=1
M1077 788 131 803 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=600 $D=1
M1078 789 131 804 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=5230 $D=1
M1079 790 131 805 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=9860 $D=1
M1080 806 800 785 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=600 $D=1
M1081 807 801 786 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=5230 $D=1
M1082 808 802 787 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=9860 $D=1
M1083 797 131 806 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=600 $D=1
M1084 798 131 807 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=5230 $D=1
M1085 799 131 808 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=9860 $D=1
M1086 809 132 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=600 $D=1
M1087 810 132 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=5230 $D=1
M1088 811 132 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=9860 $D=1
M1089 812 809 806 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=600 $D=1
M1090 813 810 807 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=5230 $D=1
M1091 814 811 808 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=9860 $D=1
M1092 803 132 812 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=600 $D=1
M1093 804 132 813 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=5230 $D=1
M1094 805 132 814 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=9860 $D=1
M1095 17 812 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=600 $D=1
M1096 18 813 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=5230 $D=1
M1097 19 814 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=9860 $D=1
M1098 815 133 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=600 $D=1
M1099 816 133 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=5230 $D=1
M1100 817 133 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=9860 $D=1
M1101 818 815 134 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=600 $D=1
M1102 819 816 135 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=5230 $D=1
M1103 820 817 136 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=9860 $D=1
M1104 137 133 818 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=600 $D=1
M1105 138 133 819 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=5230 $D=1
M1106 134 133 820 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=9860 $D=1
M1107 821 133 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=600 $D=1
M1108 822 133 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=5230 $D=1
M1109 823 133 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=9860 $D=1
M1110 830 821 139 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=600 $D=1
M1111 831 822 140 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=5230 $D=1
M1112 832 823 141 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=9860 $D=1
M1113 137 133 830 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=600 $D=1
M1114 137 133 831 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=5230 $D=1
M1115 142 133 832 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=9860 $D=1
M1116 833 133 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=600 $D=1
M1117 834 133 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=5230 $D=1
M1118 835 133 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=9860 $D=1
M1119 836 833 130 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=600 $D=1
M1120 837 834 129 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=5230 $D=1
M1121 838 835 128 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=9860 $D=1
M1122 137 133 836 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=600 $D=1
M1123 137 133 837 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=5230 $D=1
M1124 137 133 838 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=9860 $D=1
M1125 839 133 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=600 $D=1
M1126 840 133 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=5230 $D=1
M1127 841 133 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=9860 $D=1
M1128 842 839 143 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=600 $D=1
M1129 843 840 144 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=5230 $D=1
M1130 844 841 145 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=9860 $D=1
M1131 137 133 842 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=600 $D=1
M1132 137 133 843 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=5230 $D=1
M1133 137 133 844 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=9860 $D=1
M1134 845 133 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=600 $D=1
M1135 846 133 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=5230 $D=1
M1136 847 133 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=9860 $D=1
M1137 848 845 146 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=600 $D=1
M1138 849 846 147 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=5230 $D=1
M1139 850 847 148 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=9860 $D=1
M1140 137 133 848 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=600 $D=1
M1141 137 133 849 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=5230 $D=1
M1142 137 133 850 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=9860 $D=1
M1143 7 737 1080 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=600 $D=1
M1144 8 738 1081 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=5230 $D=1
M1145 9 739 1082 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=9860 $D=1
M1146 138 1080 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=600 $D=1
M1147 134 1081 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=5230 $D=1
M1148 135 1082 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=9860 $D=1
M1149 851 149 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=600 $D=1
M1150 852 149 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=5230 $D=1
M1151 853 149 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=9860 $D=1
M1152 150 851 138 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=600 $D=1
M1153 151 852 134 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=5230 $D=1
M1154 139 853 135 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=9860 $D=1
M1155 818 149 150 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=600 $D=1
M1156 819 149 151 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=5230 $D=1
M1157 820 149 139 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=9860 $D=1
M1158 854 152 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=600 $D=1
M1159 855 152 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=5230 $D=1
M1160 856 152 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=9860 $D=1
M1161 153 854 150 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=600 $D=1
M1162 154 855 151 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=5230 $D=1
M1163 155 856 139 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=9860 $D=1
M1164 830 152 153 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=600 $D=1
M1165 831 152 154 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=5230 $D=1
M1166 832 152 155 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=9860 $D=1
M1167 857 156 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=600 $D=1
M1168 858 156 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=5230 $D=1
M1169 859 156 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=9860 $D=1
M1170 157 857 153 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=600 $D=1
M1171 158 858 154 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=5230 $D=1
M1172 159 859 155 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=9860 $D=1
M1173 836 156 157 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=600 $D=1
M1174 837 156 158 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=5230 $D=1
M1175 838 156 159 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=9860 $D=1
M1176 860 160 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=600 $D=1
M1177 861 160 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=5230 $D=1
M1178 862 160 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=9860 $D=1
M1179 161 860 157 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=600 $D=1
M1180 162 861 158 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=5230 $D=1
M1181 163 862 159 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=9860 $D=1
M1182 842 160 161 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=600 $D=1
M1183 843 160 162 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=5230 $D=1
M1184 844 160 163 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=9860 $D=1
M1185 863 164 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=600 $D=1
M1186 864 164 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=5230 $D=1
M1187 865 164 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=9860 $D=1
M1188 213 863 161 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=600 $D=1
M1189 214 864 162 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=5230 $D=1
M1190 215 865 163 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=9860 $D=1
M1191 848 164 213 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=600 $D=1
M1192 849 164 214 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=5230 $D=1
M1193 850 164 215 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=9860 $D=1
M1194 866 165 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=600 $D=1
M1195 867 165 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=5230 $D=1
M1196 868 165 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=9860 $D=1
M1197 166 866 119 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=600 $D=1
M1198 869 867 120 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=5230 $D=1
M1199 870 868 121 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=9860 $D=1
M1200 14 165 166 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=600 $D=1
M1201 15 165 869 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=5230 $D=1
M1202 16 165 870 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=9860 $D=1
M1203 1113 118 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=600 $D=1
M1204 1114 723 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=5230 $D=1
M1205 1115 724 9 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=9860 $D=1
M1206 871 166 1113 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=600 $D=1
M1207 872 869 1114 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=5230 $D=1
M1208 873 870 1115 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=9860 $D=1
M1209 877 118 874 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=600 $D=1
M1210 878 723 875 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=5230 $D=1
M1211 879 724 876 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=9860 $D=1
M1212 874 166 877 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=600 $D=1
M1213 875 869 878 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=5230 $D=1
M1214 876 870 879 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=9860 $D=1
M1215 7 871 874 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=600 $D=1
M1216 8 872 875 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=5230 $D=1
M1217 9 873 876 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=9860 $D=1
M1218 1116 167 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=600 $D=1
M1219 1117 880 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=5230 $D=1
M1220 1118 881 9 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=9860 $D=1
M1221 1083 877 1116 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=600 $D=1
M1222 1084 878 1117 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=5230 $D=1
M1223 1085 879 1118 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=9860 $D=1
M1224 880 1083 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=600 $D=1
M1225 881 1084 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=5230 $D=1
M1226 168 1085 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=9860 $D=1
M1227 882 118 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=600 $D=1
M1228 883 723 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=5230 $D=1
M1229 884 724 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=9860 $D=1
M1230 7 885 882 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=600 $D=1
M1231 8 886 883 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=5230 $D=1
M1232 9 887 884 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=9860 $D=1
M1233 885 166 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=600 $D=1
M1234 886 869 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=5230 $D=1
M1235 887 870 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=9860 $D=1
M1236 1119 882 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=600 $D=1
M1237 1120 883 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=5230 $D=1
M1238 1121 884 9 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=9860 $D=1
M1239 888 167 1119 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=600 $D=1
M1240 889 880 1120 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=5230 $D=1
M1241 890 881 1121 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=9860 $D=1
M1242 893 7 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=600 $D=1
M1243 894 891 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=5230 $D=1
M1244 895 892 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=9860 $D=1
M1245 1122 888 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=600 $D=1
M1246 1123 889 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=5230 $D=1
M1247 1124 890 9 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=9860 $D=1
M1248 891 893 1122 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=600 $D=1
M1249 892 894 1123 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=5230 $D=1
M1250 169 895 1124 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=9860 $D=1
M1251 898 896 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=600 $D=1
M1252 899 897 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=5230 $D=1
M1253 900 170 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=9860 $D=1
M1254 7 904 901 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=600 $D=1
M1255 8 905 902 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=5230 $D=1
M1256 9 906 903 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=9860 $D=1
M1257 907 123 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=600 $D=1
M1258 908 124 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=5230 $D=1
M1259 909 125 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=9860 $D=1
M1260 904 907 896 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=600 $D=1
M1261 905 908 897 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=5230 $D=1
M1262 906 909 170 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=9860 $D=1
M1263 898 123 904 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=600 $D=1
M1264 899 124 905 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=5230 $D=1
M1265 900 125 906 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=9860 $D=1
M1266 910 901 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=600 $D=1
M1267 911 902 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=5230 $D=1
M1268 912 903 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=9860 $D=1
M1269 913 910 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=600 $D=1
M1270 896 911 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=5230 $D=1
M1271 897 912 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=9860 $D=1
M1272 123 901 913 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=600 $D=1
M1273 124 902 896 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=5230 $D=1
M1274 125 903 897 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=9860 $D=1
M1275 914 913 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=600 $D=1
M1276 915 896 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=5230 $D=1
M1277 916 897 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=9860 $D=1
M1278 917 901 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=600 $D=1
M1279 918 902 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=5230 $D=1
M1280 919 903 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=9860 $D=1
M1281 216 917 914 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=600 $D=1
M1282 217 918 915 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=5230 $D=1
M1283 218 919 916 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=9860 $D=1
M1284 7 901 216 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=600 $D=1
M1285 8 902 217 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=5230 $D=1
M1286 9 903 218 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=9860 $D=1
M1287 920 171 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=600 $D=1
M1288 921 171 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=5230 $D=1
M1289 922 171 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=9860 $D=1
M1290 923 920 216 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=600 $D=1
M1291 924 921 217 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=5230 $D=1
M1292 925 922 218 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=9860 $D=1
M1293 17 171 923 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=600 $D=1
M1294 18 171 924 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=5230 $D=1
M1295 19 171 925 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=9860 $D=1
M1296 926 172 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=600 $D=1
M1297 927 172 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=5230 $D=1
M1298 928 172 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=9860 $D=1
M1299 929 926 923 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=600 $D=1
M1300 172 927 924 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=5230 $D=1
M1301 172 928 925 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=9860 $D=1
M1302 7 172 929 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=600 $D=1
M1303 173 172 172 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=5230 $D=1
M1304 174 172 172 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=9860 $D=1
M1305 930 117 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=600 $D=1
M1306 931 117 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=5230 $D=1
M1307 932 117 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=9860 $D=1
M1308 7 930 933 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=600 $D=1
M1309 8 931 934 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=5230 $D=1
M1310 9 932 935 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=9860 $D=1
M1311 936 117 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=600 $D=1
M1312 937 117 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=5230 $D=1
M1313 938 117 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=9860 $D=1
M1314 939 930 929 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=600 $D=1
M1315 940 931 172 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=5230 $D=1
M1316 941 932 172 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=9860 $D=1
M1317 7 939 1086 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=600 $D=1
M1318 8 940 1087 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=5230 $D=1
M1319 9 941 1088 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=9860 $D=1
M1320 942 1086 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=600 $D=1
M1321 943 1087 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=5230 $D=1
M1322 944 1088 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=9860 $D=1
M1323 939 933 942 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=600 $D=1
M1324 940 934 943 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=5230 $D=1
M1325 941 935 944 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=9860 $D=1
M1326 945 117 942 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=600 $D=1
M1327 946 117 943 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=5230 $D=1
M1328 947 117 944 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=9860 $D=1
M1329 7 951 948 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=600 $D=1
M1330 8 952 949 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=5230 $D=1
M1331 9 953 950 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=9860 $D=1
M1332 951 117 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=600 $D=1
M1333 952 117 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=5230 $D=1
M1334 953 117 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=9860 $D=1
M1335 1089 945 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=600 $D=1
M1336 1090 946 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=5230 $D=1
M1337 1091 947 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=9860 $D=1
M1338 954 948 1089 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=600 $D=1
M1339 955 949 1090 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=5230 $D=1
M1340 956 950 1091 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=9860 $D=1
M1341 7 954 123 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=600 $D=1
M1342 8 955 124 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=5230 $D=1
M1343 9 956 125 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=9860 $D=1
M1344 1092 123 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=600 $D=1
M1345 1093 124 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=5230 $D=1
M1346 1094 125 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=9860 $D=1
M1347 954 951 1092 7 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=600 $D=1
M1348 955 952 1093 8 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=5230 $D=1
M1349 956 953 1094 9 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=9860 $D=1
M1350 177 1 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=1850 $D=0
M1351 178 1 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=6480 $D=0
M1352 179 1 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=11110 $D=0
M1353 180 1 2 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=1850 $D=0
M1354 181 1 3 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=6480 $D=0
M1355 182 1 4 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=11110 $D=0
M1356 7 177 180 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=1850 $D=0
M1357 8 178 181 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=6480 $D=0
M1358 9 179 182 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=11110 $D=0
M1359 183 1 5 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=1850 $D=0
M1360 184 1 5 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=6480 $D=0
M1361 185 1 5 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=11110 $D=0
M1362 6 177 183 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=1850 $D=0
M1363 6 178 184 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=6480 $D=0
M1364 6 179 185 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=11110 $D=0
M1365 186 1 7 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=1850 $D=0
M1366 187 1 8 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=6480 $D=0
M1367 188 1 9 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=11110 $D=0
M1368 7 177 186 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=1850 $D=0
M1369 8 178 187 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=6480 $D=0
M1370 9 179 188 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=11110 $D=0
M1371 192 11 186 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=1850 $D=0
M1372 193 11 187 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=6480 $D=0
M1373 194 11 188 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=11110 $D=0
M1374 189 11 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=1850 $D=0
M1375 190 11 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=6480 $D=0
M1376 191 11 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=11110 $D=0
M1377 195 11 183 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=1850 $D=0
M1378 196 11 184 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=6480 $D=0
M1379 197 11 185 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=11110 $D=0
M1380 180 189 195 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=1850 $D=0
M1381 181 190 196 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=6480 $D=0
M1382 182 191 197 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=11110 $D=0
M1383 198 12 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=1850 $D=0
M1384 199 12 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=6480 $D=0
M1385 200 12 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=11110 $D=0
M1386 201 12 195 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=1850 $D=0
M1387 202 12 196 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=6480 $D=0
M1388 203 12 197 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=11110 $D=0
M1389 192 198 201 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=1850 $D=0
M1390 193 199 202 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=6480 $D=0
M1391 194 200 203 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=11110 $D=0
M1392 204 13 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=1850 $D=0
M1393 205 13 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=6480 $D=0
M1394 206 13 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=11110 $D=0
M1395 207 13 7 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=1850 $D=0
M1396 208 13 8 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=6480 $D=0
M1397 209 13 9 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=11110 $D=0
M1398 14 204 207 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=1850 $D=0
M1399 15 205 208 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=6480 $D=0
M1400 16 206 209 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=11110 $D=0
M1401 210 13 17 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=1850 $D=0
M1402 211 13 18 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=6480 $D=0
M1403 212 13 19 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=11110 $D=0
M1404 213 204 210 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=1850 $D=0
M1405 214 205 211 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=6480 $D=0
M1406 215 206 212 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=11110 $D=0
M1407 219 13 216 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=1850 $D=0
M1408 220 13 217 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=6480 $D=0
M1409 221 13 218 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=11110 $D=0
M1410 201 204 219 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=1850 $D=0
M1411 202 205 220 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=6480 $D=0
M1412 203 206 221 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=11110 $D=0
M1413 225 20 219 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=1850 $D=0
M1414 226 20 220 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=6480 $D=0
M1415 227 20 221 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=11110 $D=0
M1416 222 20 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=1850 $D=0
M1417 223 20 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=6480 $D=0
M1418 224 20 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=11110 $D=0
M1419 228 20 210 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=1850 $D=0
M1420 229 20 211 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=6480 $D=0
M1421 230 20 212 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=11110 $D=0
M1422 207 222 228 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=1850 $D=0
M1423 208 223 229 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=6480 $D=0
M1424 209 224 230 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=11110 $D=0
M1425 231 21 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=1850 $D=0
M1426 232 21 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=6480 $D=0
M1427 233 21 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=11110 $D=0
M1428 234 21 228 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=1850 $D=0
M1429 235 21 229 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=6480 $D=0
M1430 236 21 230 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=11110 $D=0
M1431 225 231 234 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=1850 $D=0
M1432 226 232 235 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=6480 $D=0
M1433 227 233 236 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=11110 $D=0
M1434 167 22 237 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=1850 $D=0
M1435 173 22 238 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=6480 $D=0
M1436 174 22 239 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=11110 $D=0
M1437 240 23 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=1850 $D=0
M1438 241 23 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=6480 $D=0
M1439 242 23 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=11110 $D=0
M1440 243 237 234 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=1850 $D=0
M1441 244 238 235 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=6480 $D=0
M1442 245 239 236 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=11110 $D=0
M1443 167 243 957 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=1850 $D=0
M1444 173 244 958 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=6480 $D=0
M1445 174 245 959 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=11110 $D=0
M1446 246 957 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=1850 $D=0
M1447 247 958 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=6480 $D=0
M1448 248 959 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=11110 $D=0
M1449 243 22 246 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=1850 $D=0
M1450 244 22 247 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=6480 $D=0
M1451 245 22 248 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=11110 $D=0
M1452 246 240 249 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=1850 $D=0
M1453 247 241 250 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=6480 $D=0
M1454 248 242 251 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=11110 $D=0
M1455 255 252 246 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=1850 $D=0
M1456 256 253 247 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=6480 $D=0
M1457 257 254 248 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=11110 $D=0
M1458 252 24 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=1850 $D=0
M1459 253 24 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=6480 $D=0
M1460 254 24 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=11110 $D=0
M1461 167 25 258 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=1850 $D=0
M1462 173 25 259 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=6480 $D=0
M1463 174 25 260 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=11110 $D=0
M1464 261 26 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=1850 $D=0
M1465 262 26 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=6480 $D=0
M1466 263 26 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=11110 $D=0
M1467 264 258 234 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=1850 $D=0
M1468 265 259 235 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=6480 $D=0
M1469 266 260 236 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=11110 $D=0
M1470 167 264 960 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=1850 $D=0
M1471 173 265 961 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=6480 $D=0
M1472 174 266 962 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=11110 $D=0
M1473 267 960 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=1850 $D=0
M1474 268 961 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=6480 $D=0
M1475 269 962 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=11110 $D=0
M1476 264 25 267 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=1850 $D=0
M1477 265 25 268 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=6480 $D=0
M1478 266 25 269 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=11110 $D=0
M1479 267 261 249 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=1850 $D=0
M1480 268 262 250 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=6480 $D=0
M1481 269 263 251 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=11110 $D=0
M1482 255 270 267 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=1850 $D=0
M1483 256 271 268 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=6480 $D=0
M1484 257 272 269 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=11110 $D=0
M1485 270 27 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=1850 $D=0
M1486 271 27 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=6480 $D=0
M1487 272 27 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=11110 $D=0
M1488 167 28 273 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=1850 $D=0
M1489 173 28 274 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=6480 $D=0
M1490 174 28 275 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=11110 $D=0
M1491 276 29 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=1850 $D=0
M1492 277 29 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=6480 $D=0
M1493 278 29 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=11110 $D=0
M1494 279 273 234 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=1850 $D=0
M1495 280 274 235 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=6480 $D=0
M1496 281 275 236 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=11110 $D=0
M1497 167 279 963 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=1850 $D=0
M1498 173 280 964 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=6480 $D=0
M1499 174 281 965 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=11110 $D=0
M1500 282 963 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=1850 $D=0
M1501 283 964 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=6480 $D=0
M1502 284 965 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=11110 $D=0
M1503 279 28 282 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=1850 $D=0
M1504 280 28 283 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=6480 $D=0
M1505 281 28 284 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=11110 $D=0
M1506 282 276 249 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=1850 $D=0
M1507 283 277 250 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=6480 $D=0
M1508 284 278 251 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=11110 $D=0
M1509 255 285 282 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=1850 $D=0
M1510 256 286 283 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=6480 $D=0
M1511 257 287 284 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=11110 $D=0
M1512 285 30 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=1850 $D=0
M1513 286 30 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=6480 $D=0
M1514 287 30 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=11110 $D=0
M1515 167 31 288 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=1850 $D=0
M1516 173 31 289 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=6480 $D=0
M1517 174 31 290 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=11110 $D=0
M1518 291 32 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=1850 $D=0
M1519 292 32 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=6480 $D=0
M1520 293 32 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=11110 $D=0
M1521 294 288 234 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=1850 $D=0
M1522 295 289 235 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=6480 $D=0
M1523 296 290 236 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=11110 $D=0
M1524 167 294 966 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=1850 $D=0
M1525 173 295 967 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=6480 $D=0
M1526 174 296 968 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=11110 $D=0
M1527 297 966 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=1850 $D=0
M1528 298 967 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=6480 $D=0
M1529 299 968 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=11110 $D=0
M1530 294 31 297 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=1850 $D=0
M1531 295 31 298 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=6480 $D=0
M1532 296 31 299 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=11110 $D=0
M1533 297 291 249 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=1850 $D=0
M1534 298 292 250 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=6480 $D=0
M1535 299 293 251 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=11110 $D=0
M1536 255 300 297 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=1850 $D=0
M1537 256 301 298 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=6480 $D=0
M1538 257 302 299 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=11110 $D=0
M1539 300 33 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=1850 $D=0
M1540 301 33 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=6480 $D=0
M1541 302 33 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=11110 $D=0
M1542 167 34 303 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=1850 $D=0
M1543 173 34 304 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=6480 $D=0
M1544 174 34 305 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=11110 $D=0
M1545 306 35 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=1850 $D=0
M1546 307 35 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=6480 $D=0
M1547 308 35 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=11110 $D=0
M1548 309 303 234 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=1850 $D=0
M1549 310 304 235 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=6480 $D=0
M1550 311 305 236 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=11110 $D=0
M1551 167 309 969 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=1850 $D=0
M1552 173 310 970 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=6480 $D=0
M1553 174 311 971 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=11110 $D=0
M1554 312 969 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=1850 $D=0
M1555 313 970 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=6480 $D=0
M1556 314 971 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=11110 $D=0
M1557 309 34 312 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=1850 $D=0
M1558 310 34 313 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=6480 $D=0
M1559 311 34 314 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=11110 $D=0
M1560 312 306 249 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=1850 $D=0
M1561 313 307 250 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=6480 $D=0
M1562 314 308 251 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=11110 $D=0
M1563 255 315 312 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=1850 $D=0
M1564 256 316 313 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=6480 $D=0
M1565 257 317 314 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=11110 $D=0
M1566 315 36 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=1850 $D=0
M1567 316 36 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=6480 $D=0
M1568 317 36 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=11110 $D=0
M1569 167 37 318 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=1850 $D=0
M1570 173 37 319 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=6480 $D=0
M1571 174 37 320 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=11110 $D=0
M1572 321 38 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=1850 $D=0
M1573 322 38 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=6480 $D=0
M1574 323 38 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=11110 $D=0
M1575 324 318 234 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=1850 $D=0
M1576 325 319 235 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=6480 $D=0
M1577 326 320 236 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=11110 $D=0
M1578 167 324 972 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=1850 $D=0
M1579 173 325 973 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=6480 $D=0
M1580 174 326 974 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=11110 $D=0
M1581 327 972 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=1850 $D=0
M1582 328 973 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=6480 $D=0
M1583 329 974 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=11110 $D=0
M1584 324 37 327 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=1850 $D=0
M1585 325 37 328 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=6480 $D=0
M1586 326 37 329 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=11110 $D=0
M1587 327 321 249 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=1850 $D=0
M1588 328 322 250 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=6480 $D=0
M1589 329 323 251 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=11110 $D=0
M1590 255 330 327 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=1850 $D=0
M1591 256 331 328 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=6480 $D=0
M1592 257 332 329 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=11110 $D=0
M1593 330 39 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=1850 $D=0
M1594 331 39 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=6480 $D=0
M1595 332 39 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=11110 $D=0
M1596 167 40 333 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=1850 $D=0
M1597 173 40 334 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=6480 $D=0
M1598 174 40 335 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=11110 $D=0
M1599 336 41 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=1850 $D=0
M1600 337 41 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=6480 $D=0
M1601 338 41 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=11110 $D=0
M1602 339 333 234 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=1850 $D=0
M1603 340 334 235 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=6480 $D=0
M1604 341 335 236 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=11110 $D=0
M1605 167 339 975 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=1850 $D=0
M1606 173 340 976 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=6480 $D=0
M1607 174 341 977 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=11110 $D=0
M1608 342 975 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=1850 $D=0
M1609 343 976 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=6480 $D=0
M1610 344 977 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=11110 $D=0
M1611 339 40 342 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=1850 $D=0
M1612 340 40 343 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=6480 $D=0
M1613 341 40 344 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=11110 $D=0
M1614 342 336 249 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=1850 $D=0
M1615 343 337 250 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=6480 $D=0
M1616 344 338 251 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=11110 $D=0
M1617 255 345 342 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=1850 $D=0
M1618 256 346 343 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=6480 $D=0
M1619 257 347 344 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=11110 $D=0
M1620 345 42 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=1850 $D=0
M1621 346 42 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=6480 $D=0
M1622 347 42 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=11110 $D=0
M1623 167 43 348 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=1850 $D=0
M1624 173 43 349 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=6480 $D=0
M1625 174 43 350 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=11110 $D=0
M1626 351 44 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=1850 $D=0
M1627 352 44 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=6480 $D=0
M1628 353 44 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=11110 $D=0
M1629 354 348 234 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=1850 $D=0
M1630 355 349 235 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=6480 $D=0
M1631 356 350 236 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=11110 $D=0
M1632 167 354 978 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=1850 $D=0
M1633 173 355 979 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=6480 $D=0
M1634 174 356 980 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=11110 $D=0
M1635 357 978 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=1850 $D=0
M1636 358 979 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=6480 $D=0
M1637 359 980 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=11110 $D=0
M1638 354 43 357 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=1850 $D=0
M1639 355 43 358 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=6480 $D=0
M1640 356 43 359 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=11110 $D=0
M1641 357 351 249 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=1850 $D=0
M1642 358 352 250 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=6480 $D=0
M1643 359 353 251 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=11110 $D=0
M1644 255 360 357 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=1850 $D=0
M1645 256 361 358 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=6480 $D=0
M1646 257 362 359 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=11110 $D=0
M1647 360 45 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=1850 $D=0
M1648 361 45 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=6480 $D=0
M1649 362 45 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=11110 $D=0
M1650 167 46 363 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=1850 $D=0
M1651 173 46 364 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=6480 $D=0
M1652 174 46 365 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=11110 $D=0
M1653 366 47 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=1850 $D=0
M1654 367 47 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=6480 $D=0
M1655 368 47 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=11110 $D=0
M1656 369 363 234 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=1850 $D=0
M1657 370 364 235 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=6480 $D=0
M1658 371 365 236 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=11110 $D=0
M1659 167 369 981 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=1850 $D=0
M1660 173 370 982 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=6480 $D=0
M1661 174 371 983 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=11110 $D=0
M1662 372 981 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=1850 $D=0
M1663 373 982 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=6480 $D=0
M1664 374 983 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=11110 $D=0
M1665 369 46 372 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=1850 $D=0
M1666 370 46 373 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=6480 $D=0
M1667 371 46 374 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=11110 $D=0
M1668 372 366 249 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=1850 $D=0
M1669 373 367 250 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=6480 $D=0
M1670 374 368 251 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=11110 $D=0
M1671 255 375 372 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=1850 $D=0
M1672 256 376 373 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=6480 $D=0
M1673 257 377 374 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=11110 $D=0
M1674 375 48 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=1850 $D=0
M1675 376 48 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=6480 $D=0
M1676 377 48 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=11110 $D=0
M1677 167 49 378 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=1850 $D=0
M1678 173 49 379 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=6480 $D=0
M1679 174 49 380 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=11110 $D=0
M1680 381 50 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=1850 $D=0
M1681 382 50 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=6480 $D=0
M1682 383 50 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=11110 $D=0
M1683 384 378 234 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=1850 $D=0
M1684 385 379 235 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=6480 $D=0
M1685 386 380 236 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=11110 $D=0
M1686 167 384 984 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=1850 $D=0
M1687 173 385 985 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=6480 $D=0
M1688 174 386 986 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=11110 $D=0
M1689 387 984 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=1850 $D=0
M1690 388 985 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=6480 $D=0
M1691 389 986 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=11110 $D=0
M1692 384 49 387 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=1850 $D=0
M1693 385 49 388 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=6480 $D=0
M1694 386 49 389 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=11110 $D=0
M1695 387 381 249 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=1850 $D=0
M1696 388 382 250 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=6480 $D=0
M1697 389 383 251 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=11110 $D=0
M1698 255 390 387 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=1850 $D=0
M1699 256 391 388 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=6480 $D=0
M1700 257 392 389 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=11110 $D=0
M1701 390 51 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=1850 $D=0
M1702 391 51 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=6480 $D=0
M1703 392 51 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=11110 $D=0
M1704 167 52 393 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=1850 $D=0
M1705 173 52 394 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=6480 $D=0
M1706 174 52 395 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=11110 $D=0
M1707 396 53 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=1850 $D=0
M1708 397 53 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=6480 $D=0
M1709 398 53 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=11110 $D=0
M1710 399 393 234 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=1850 $D=0
M1711 400 394 235 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=6480 $D=0
M1712 401 395 236 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=11110 $D=0
M1713 167 399 987 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=1850 $D=0
M1714 173 400 988 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=6480 $D=0
M1715 174 401 989 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=11110 $D=0
M1716 402 987 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=1850 $D=0
M1717 403 988 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=6480 $D=0
M1718 404 989 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=11110 $D=0
M1719 399 52 402 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=1850 $D=0
M1720 400 52 403 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=6480 $D=0
M1721 401 52 404 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=11110 $D=0
M1722 402 396 249 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=1850 $D=0
M1723 403 397 250 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=6480 $D=0
M1724 404 398 251 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=11110 $D=0
M1725 255 405 402 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=1850 $D=0
M1726 256 406 403 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=6480 $D=0
M1727 257 407 404 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=11110 $D=0
M1728 405 54 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=1850 $D=0
M1729 406 54 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=6480 $D=0
M1730 407 54 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=11110 $D=0
M1731 167 55 408 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=1850 $D=0
M1732 173 55 409 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=6480 $D=0
M1733 174 55 410 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=11110 $D=0
M1734 411 56 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=1850 $D=0
M1735 412 56 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=6480 $D=0
M1736 413 56 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=11110 $D=0
M1737 414 408 234 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=1850 $D=0
M1738 415 409 235 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=6480 $D=0
M1739 416 410 236 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=11110 $D=0
M1740 167 414 990 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=1850 $D=0
M1741 173 415 991 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=6480 $D=0
M1742 174 416 992 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=11110 $D=0
M1743 417 990 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=1850 $D=0
M1744 418 991 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=6480 $D=0
M1745 419 992 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=11110 $D=0
M1746 414 55 417 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=1850 $D=0
M1747 415 55 418 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=6480 $D=0
M1748 416 55 419 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=11110 $D=0
M1749 417 411 249 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=1850 $D=0
M1750 418 412 250 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=6480 $D=0
M1751 419 413 251 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=11110 $D=0
M1752 255 420 417 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=1850 $D=0
M1753 256 421 418 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=6480 $D=0
M1754 257 422 419 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=11110 $D=0
M1755 420 57 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=1850 $D=0
M1756 421 57 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=6480 $D=0
M1757 422 57 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=11110 $D=0
M1758 167 58 423 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=1850 $D=0
M1759 173 58 424 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=6480 $D=0
M1760 174 58 425 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=11110 $D=0
M1761 426 59 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=1850 $D=0
M1762 427 59 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=6480 $D=0
M1763 428 59 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=11110 $D=0
M1764 429 423 234 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=1850 $D=0
M1765 430 424 235 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=6480 $D=0
M1766 431 425 236 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=11110 $D=0
M1767 167 429 993 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=1850 $D=0
M1768 173 430 994 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=6480 $D=0
M1769 174 431 995 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=11110 $D=0
M1770 432 993 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=1850 $D=0
M1771 433 994 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=6480 $D=0
M1772 434 995 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=11110 $D=0
M1773 429 58 432 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=1850 $D=0
M1774 430 58 433 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=6480 $D=0
M1775 431 58 434 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=11110 $D=0
M1776 432 426 249 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=1850 $D=0
M1777 433 427 250 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=6480 $D=0
M1778 434 428 251 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=11110 $D=0
M1779 255 435 432 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=1850 $D=0
M1780 256 436 433 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=6480 $D=0
M1781 257 437 434 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=11110 $D=0
M1782 435 60 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=1850 $D=0
M1783 436 60 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=6480 $D=0
M1784 437 60 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=11110 $D=0
M1785 167 61 438 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=1850 $D=0
M1786 173 61 439 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=6480 $D=0
M1787 174 61 440 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=11110 $D=0
M1788 441 62 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=1850 $D=0
M1789 442 62 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=6480 $D=0
M1790 443 62 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=11110 $D=0
M1791 444 438 234 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=1850 $D=0
M1792 445 439 235 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=6480 $D=0
M1793 446 440 236 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=11110 $D=0
M1794 167 444 996 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=1850 $D=0
M1795 173 445 997 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=6480 $D=0
M1796 174 446 998 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=11110 $D=0
M1797 447 996 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=1850 $D=0
M1798 448 997 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=6480 $D=0
M1799 449 998 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=11110 $D=0
M1800 444 61 447 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=1850 $D=0
M1801 445 61 448 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=6480 $D=0
M1802 446 61 449 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=11110 $D=0
M1803 447 441 249 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=1850 $D=0
M1804 448 442 250 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=6480 $D=0
M1805 449 443 251 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=11110 $D=0
M1806 255 450 447 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=1850 $D=0
M1807 256 451 448 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=6480 $D=0
M1808 257 452 449 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=11110 $D=0
M1809 450 63 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=1850 $D=0
M1810 451 63 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=6480 $D=0
M1811 452 63 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=11110 $D=0
M1812 167 64 453 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=1850 $D=0
M1813 173 64 454 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=6480 $D=0
M1814 174 64 455 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=11110 $D=0
M1815 456 65 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=1850 $D=0
M1816 457 65 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=6480 $D=0
M1817 458 65 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=11110 $D=0
M1818 459 453 234 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=1850 $D=0
M1819 460 454 235 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=6480 $D=0
M1820 461 455 236 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=11110 $D=0
M1821 167 459 999 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=1850 $D=0
M1822 173 460 1000 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=6480 $D=0
M1823 174 461 1001 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=11110 $D=0
M1824 462 999 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=1850 $D=0
M1825 463 1000 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=6480 $D=0
M1826 464 1001 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=11110 $D=0
M1827 459 64 462 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=1850 $D=0
M1828 460 64 463 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=6480 $D=0
M1829 461 64 464 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=11110 $D=0
M1830 462 456 249 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=1850 $D=0
M1831 463 457 250 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=6480 $D=0
M1832 464 458 251 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=11110 $D=0
M1833 255 465 462 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=1850 $D=0
M1834 256 466 463 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=6480 $D=0
M1835 257 467 464 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=11110 $D=0
M1836 465 66 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=1850 $D=0
M1837 466 66 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=6480 $D=0
M1838 467 66 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=11110 $D=0
M1839 167 67 468 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=1850 $D=0
M1840 173 67 469 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=6480 $D=0
M1841 174 67 470 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=11110 $D=0
M1842 471 68 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=1850 $D=0
M1843 472 68 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=6480 $D=0
M1844 473 68 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=11110 $D=0
M1845 474 468 234 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=1850 $D=0
M1846 475 469 235 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=6480 $D=0
M1847 476 470 236 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=11110 $D=0
M1848 167 474 1002 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=1850 $D=0
M1849 173 475 1003 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=6480 $D=0
M1850 174 476 1004 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=11110 $D=0
M1851 477 1002 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=1850 $D=0
M1852 478 1003 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=6480 $D=0
M1853 479 1004 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=11110 $D=0
M1854 474 67 477 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=1850 $D=0
M1855 475 67 478 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=6480 $D=0
M1856 476 67 479 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=11110 $D=0
M1857 477 471 249 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=1850 $D=0
M1858 478 472 250 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=6480 $D=0
M1859 479 473 251 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=11110 $D=0
M1860 255 480 477 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=1850 $D=0
M1861 256 481 478 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=6480 $D=0
M1862 257 482 479 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=11110 $D=0
M1863 480 69 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=1850 $D=0
M1864 481 69 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=6480 $D=0
M1865 482 69 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=11110 $D=0
M1866 167 70 483 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=1850 $D=0
M1867 173 70 484 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=6480 $D=0
M1868 174 70 485 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=11110 $D=0
M1869 486 71 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=1850 $D=0
M1870 487 71 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=6480 $D=0
M1871 488 71 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=11110 $D=0
M1872 489 483 234 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=1850 $D=0
M1873 490 484 235 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=6480 $D=0
M1874 491 485 236 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=11110 $D=0
M1875 167 489 1005 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=1850 $D=0
M1876 173 490 1006 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=6480 $D=0
M1877 174 491 1007 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=11110 $D=0
M1878 492 1005 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=1850 $D=0
M1879 493 1006 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=6480 $D=0
M1880 494 1007 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=11110 $D=0
M1881 489 70 492 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=1850 $D=0
M1882 490 70 493 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=6480 $D=0
M1883 491 70 494 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=11110 $D=0
M1884 492 486 249 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=1850 $D=0
M1885 493 487 250 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=6480 $D=0
M1886 494 488 251 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=11110 $D=0
M1887 255 495 492 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=1850 $D=0
M1888 256 496 493 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=6480 $D=0
M1889 257 497 494 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=11110 $D=0
M1890 495 72 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=1850 $D=0
M1891 496 72 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=6480 $D=0
M1892 497 72 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=11110 $D=0
M1893 167 73 498 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=1850 $D=0
M1894 173 73 499 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=6480 $D=0
M1895 174 73 500 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=11110 $D=0
M1896 501 74 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=1850 $D=0
M1897 502 74 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=6480 $D=0
M1898 503 74 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=11110 $D=0
M1899 504 498 234 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=1850 $D=0
M1900 505 499 235 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=6480 $D=0
M1901 506 500 236 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=11110 $D=0
M1902 167 504 1008 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=1850 $D=0
M1903 173 505 1009 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=6480 $D=0
M1904 174 506 1010 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=11110 $D=0
M1905 507 1008 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=1850 $D=0
M1906 508 1009 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=6480 $D=0
M1907 509 1010 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=11110 $D=0
M1908 504 73 507 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=1850 $D=0
M1909 505 73 508 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=6480 $D=0
M1910 506 73 509 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=11110 $D=0
M1911 507 501 249 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=1850 $D=0
M1912 508 502 250 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=6480 $D=0
M1913 509 503 251 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=11110 $D=0
M1914 255 510 507 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=1850 $D=0
M1915 256 511 508 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=6480 $D=0
M1916 257 512 509 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=11110 $D=0
M1917 510 75 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=1850 $D=0
M1918 511 75 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=6480 $D=0
M1919 512 75 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=11110 $D=0
M1920 167 76 513 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=1850 $D=0
M1921 173 76 514 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=6480 $D=0
M1922 174 76 515 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=11110 $D=0
M1923 516 77 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=1850 $D=0
M1924 517 77 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=6480 $D=0
M1925 518 77 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=11110 $D=0
M1926 519 513 234 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=1850 $D=0
M1927 520 514 235 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=6480 $D=0
M1928 521 515 236 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=11110 $D=0
M1929 167 519 1011 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=1850 $D=0
M1930 173 520 1012 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=6480 $D=0
M1931 174 521 1013 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=11110 $D=0
M1932 522 1011 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=1850 $D=0
M1933 523 1012 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=6480 $D=0
M1934 524 1013 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=11110 $D=0
M1935 519 76 522 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=1850 $D=0
M1936 520 76 523 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=6480 $D=0
M1937 521 76 524 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=11110 $D=0
M1938 522 516 249 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=1850 $D=0
M1939 523 517 250 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=6480 $D=0
M1940 524 518 251 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=11110 $D=0
M1941 255 525 522 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=1850 $D=0
M1942 256 526 523 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=6480 $D=0
M1943 257 527 524 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=11110 $D=0
M1944 525 78 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=1850 $D=0
M1945 526 78 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=6480 $D=0
M1946 527 78 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=11110 $D=0
M1947 167 79 528 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=1850 $D=0
M1948 173 79 529 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=6480 $D=0
M1949 174 79 530 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=11110 $D=0
M1950 531 80 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=1850 $D=0
M1951 532 80 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=6480 $D=0
M1952 533 80 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=11110 $D=0
M1953 534 528 234 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=1850 $D=0
M1954 535 529 235 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=6480 $D=0
M1955 536 530 236 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=11110 $D=0
M1956 167 534 1014 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=1850 $D=0
M1957 173 535 1015 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=6480 $D=0
M1958 174 536 1016 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=11110 $D=0
M1959 537 1014 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=1850 $D=0
M1960 538 1015 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=6480 $D=0
M1961 539 1016 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=11110 $D=0
M1962 534 79 537 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=1850 $D=0
M1963 535 79 538 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=6480 $D=0
M1964 536 79 539 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=11110 $D=0
M1965 537 531 249 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=1850 $D=0
M1966 538 532 250 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=6480 $D=0
M1967 539 533 251 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=11110 $D=0
M1968 255 540 537 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=1850 $D=0
M1969 256 541 538 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=6480 $D=0
M1970 257 542 539 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=11110 $D=0
M1971 540 81 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=1850 $D=0
M1972 541 81 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=6480 $D=0
M1973 542 81 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=11110 $D=0
M1974 167 82 543 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=1850 $D=0
M1975 173 82 544 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=6480 $D=0
M1976 174 82 545 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=11110 $D=0
M1977 546 83 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=1850 $D=0
M1978 547 83 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=6480 $D=0
M1979 548 83 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=11110 $D=0
M1980 549 543 234 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=1850 $D=0
M1981 550 544 235 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=6480 $D=0
M1982 551 545 236 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=11110 $D=0
M1983 167 549 1017 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=1850 $D=0
M1984 173 550 1018 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=6480 $D=0
M1985 174 551 1019 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=11110 $D=0
M1986 552 1017 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=1850 $D=0
M1987 553 1018 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=6480 $D=0
M1988 554 1019 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=11110 $D=0
M1989 549 82 552 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=1850 $D=0
M1990 550 82 553 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=6480 $D=0
M1991 551 82 554 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=11110 $D=0
M1992 552 546 249 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=1850 $D=0
M1993 553 547 250 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=6480 $D=0
M1994 554 548 251 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=11110 $D=0
M1995 255 555 552 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=1850 $D=0
M1996 256 556 553 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=6480 $D=0
M1997 257 557 554 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=11110 $D=0
M1998 555 84 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=1850 $D=0
M1999 556 84 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=6480 $D=0
M2000 557 84 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=11110 $D=0
M2001 167 85 558 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=1850 $D=0
M2002 173 85 559 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=6480 $D=0
M2003 174 85 560 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=11110 $D=0
M2004 561 86 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=1850 $D=0
M2005 562 86 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=6480 $D=0
M2006 563 86 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=11110 $D=0
M2007 564 558 234 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=1850 $D=0
M2008 565 559 235 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=6480 $D=0
M2009 566 560 236 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=11110 $D=0
M2010 167 564 1020 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=1850 $D=0
M2011 173 565 1021 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=6480 $D=0
M2012 174 566 1022 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=11110 $D=0
M2013 567 1020 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=1850 $D=0
M2014 568 1021 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=6480 $D=0
M2015 569 1022 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=11110 $D=0
M2016 564 85 567 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=1850 $D=0
M2017 565 85 568 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=6480 $D=0
M2018 566 85 569 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=11110 $D=0
M2019 567 561 249 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=1850 $D=0
M2020 568 562 250 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=6480 $D=0
M2021 569 563 251 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=11110 $D=0
M2022 255 570 567 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=1850 $D=0
M2023 256 571 568 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=6480 $D=0
M2024 257 572 569 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=11110 $D=0
M2025 570 87 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=1850 $D=0
M2026 571 87 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=6480 $D=0
M2027 572 87 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=11110 $D=0
M2028 167 88 573 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=1850 $D=0
M2029 173 88 574 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=6480 $D=0
M2030 174 88 575 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=11110 $D=0
M2031 576 89 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=1850 $D=0
M2032 577 89 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=6480 $D=0
M2033 578 89 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=11110 $D=0
M2034 579 573 234 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=1850 $D=0
M2035 580 574 235 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=6480 $D=0
M2036 581 575 236 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=11110 $D=0
M2037 167 579 1023 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=1850 $D=0
M2038 173 580 1024 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=6480 $D=0
M2039 174 581 1025 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=11110 $D=0
M2040 582 1023 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=1850 $D=0
M2041 583 1024 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=6480 $D=0
M2042 584 1025 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=11110 $D=0
M2043 579 88 582 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=1850 $D=0
M2044 580 88 583 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=6480 $D=0
M2045 581 88 584 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=11110 $D=0
M2046 582 576 249 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=1850 $D=0
M2047 583 577 250 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=6480 $D=0
M2048 584 578 251 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=11110 $D=0
M2049 255 585 582 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=1850 $D=0
M2050 256 586 583 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=6480 $D=0
M2051 257 587 584 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=11110 $D=0
M2052 585 90 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=1850 $D=0
M2053 586 90 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=6480 $D=0
M2054 587 90 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=11110 $D=0
M2055 167 91 588 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=1850 $D=0
M2056 173 91 589 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=6480 $D=0
M2057 174 91 590 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=11110 $D=0
M2058 591 92 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=1850 $D=0
M2059 592 92 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=6480 $D=0
M2060 593 92 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=11110 $D=0
M2061 594 588 234 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=1850 $D=0
M2062 595 589 235 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=6480 $D=0
M2063 596 590 236 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=11110 $D=0
M2064 167 594 1026 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=1850 $D=0
M2065 173 595 1027 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=6480 $D=0
M2066 174 596 1028 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=11110 $D=0
M2067 597 1026 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=1850 $D=0
M2068 598 1027 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=6480 $D=0
M2069 599 1028 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=11110 $D=0
M2070 594 91 597 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=1850 $D=0
M2071 595 91 598 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=6480 $D=0
M2072 596 91 599 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=11110 $D=0
M2073 597 591 249 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=1850 $D=0
M2074 598 592 250 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=6480 $D=0
M2075 599 593 251 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=11110 $D=0
M2076 255 600 597 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=1850 $D=0
M2077 256 601 598 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=6480 $D=0
M2078 257 602 599 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=11110 $D=0
M2079 600 93 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=1850 $D=0
M2080 601 93 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=6480 $D=0
M2081 602 93 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=11110 $D=0
M2082 167 94 603 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=1850 $D=0
M2083 173 94 604 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=6480 $D=0
M2084 174 94 605 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=11110 $D=0
M2085 606 95 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=1850 $D=0
M2086 607 95 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=6480 $D=0
M2087 608 95 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=11110 $D=0
M2088 609 603 234 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=1850 $D=0
M2089 610 604 235 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=6480 $D=0
M2090 611 605 236 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=11110 $D=0
M2091 167 609 1029 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=1850 $D=0
M2092 173 610 1030 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=6480 $D=0
M2093 174 611 1031 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=11110 $D=0
M2094 612 1029 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=1850 $D=0
M2095 613 1030 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=6480 $D=0
M2096 614 1031 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=11110 $D=0
M2097 609 94 612 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=1850 $D=0
M2098 610 94 613 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=6480 $D=0
M2099 611 94 614 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=11110 $D=0
M2100 612 606 249 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=1850 $D=0
M2101 613 607 250 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=6480 $D=0
M2102 614 608 251 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=11110 $D=0
M2103 255 615 612 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=1850 $D=0
M2104 256 616 613 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=6480 $D=0
M2105 257 617 614 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=11110 $D=0
M2106 615 96 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=1850 $D=0
M2107 616 96 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=6480 $D=0
M2108 617 96 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=11110 $D=0
M2109 167 97 618 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=1850 $D=0
M2110 173 97 619 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=6480 $D=0
M2111 174 97 620 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=11110 $D=0
M2112 621 98 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=1850 $D=0
M2113 622 98 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=6480 $D=0
M2114 623 98 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=11110 $D=0
M2115 624 618 234 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=1850 $D=0
M2116 625 619 235 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=6480 $D=0
M2117 626 620 236 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=11110 $D=0
M2118 167 624 1032 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=1850 $D=0
M2119 173 625 1033 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=6480 $D=0
M2120 174 626 1034 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=11110 $D=0
M2121 627 1032 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=1850 $D=0
M2122 628 1033 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=6480 $D=0
M2123 629 1034 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=11110 $D=0
M2124 624 97 627 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=1850 $D=0
M2125 625 97 628 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=6480 $D=0
M2126 626 97 629 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=11110 $D=0
M2127 627 621 249 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=1850 $D=0
M2128 628 622 250 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=6480 $D=0
M2129 629 623 251 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=11110 $D=0
M2130 255 630 627 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=1850 $D=0
M2131 256 631 628 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=6480 $D=0
M2132 257 632 629 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=11110 $D=0
M2133 630 99 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=1850 $D=0
M2134 631 99 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=6480 $D=0
M2135 632 99 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=11110 $D=0
M2136 167 100 633 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=1850 $D=0
M2137 173 100 634 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=6480 $D=0
M2138 174 100 635 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=11110 $D=0
M2139 636 101 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=1850 $D=0
M2140 637 101 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=6480 $D=0
M2141 638 101 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=11110 $D=0
M2142 639 633 234 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=1850 $D=0
M2143 640 634 235 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=6480 $D=0
M2144 641 635 236 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=11110 $D=0
M2145 167 639 1035 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=1850 $D=0
M2146 173 640 1036 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=6480 $D=0
M2147 174 641 1037 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=11110 $D=0
M2148 642 1035 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=1850 $D=0
M2149 643 1036 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=6480 $D=0
M2150 644 1037 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=11110 $D=0
M2151 639 100 642 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=1850 $D=0
M2152 640 100 643 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=6480 $D=0
M2153 641 100 644 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=11110 $D=0
M2154 642 636 249 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=1850 $D=0
M2155 643 637 250 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=6480 $D=0
M2156 644 638 251 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=11110 $D=0
M2157 255 645 642 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=1850 $D=0
M2158 256 646 643 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=6480 $D=0
M2159 257 647 644 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=11110 $D=0
M2160 645 102 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=1850 $D=0
M2161 646 102 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=6480 $D=0
M2162 647 102 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=11110 $D=0
M2163 167 103 648 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=1850 $D=0
M2164 173 103 649 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=6480 $D=0
M2165 174 103 650 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=11110 $D=0
M2166 651 104 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=1850 $D=0
M2167 652 104 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=6480 $D=0
M2168 653 104 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=11110 $D=0
M2169 654 648 234 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=1850 $D=0
M2170 655 649 235 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=6480 $D=0
M2171 656 650 236 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=11110 $D=0
M2172 167 654 1038 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=1850 $D=0
M2173 173 655 1039 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=6480 $D=0
M2174 174 656 1040 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=11110 $D=0
M2175 657 1038 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=1850 $D=0
M2176 658 1039 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=6480 $D=0
M2177 659 1040 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=11110 $D=0
M2178 654 103 657 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=1850 $D=0
M2179 655 103 658 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=6480 $D=0
M2180 656 103 659 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=11110 $D=0
M2181 657 651 249 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=1850 $D=0
M2182 658 652 250 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=6480 $D=0
M2183 659 653 251 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=11110 $D=0
M2184 255 660 657 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=1850 $D=0
M2185 256 661 658 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=6480 $D=0
M2186 257 662 659 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=11110 $D=0
M2187 660 105 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=1850 $D=0
M2188 661 105 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=6480 $D=0
M2189 662 105 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=11110 $D=0
M2190 167 106 663 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=1850 $D=0
M2191 173 106 664 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=6480 $D=0
M2192 174 106 665 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=11110 $D=0
M2193 666 107 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=1850 $D=0
M2194 667 107 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=6480 $D=0
M2195 668 107 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=11110 $D=0
M2196 669 663 234 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=1850 $D=0
M2197 670 664 235 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=6480 $D=0
M2198 671 665 236 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=11110 $D=0
M2199 167 669 1041 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=1850 $D=0
M2200 173 670 1042 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=6480 $D=0
M2201 174 671 1043 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=11110 $D=0
M2202 672 1041 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=1850 $D=0
M2203 673 1042 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=6480 $D=0
M2204 674 1043 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=11110 $D=0
M2205 669 106 672 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=1850 $D=0
M2206 670 106 673 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=6480 $D=0
M2207 671 106 674 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=11110 $D=0
M2208 672 666 249 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=1850 $D=0
M2209 673 667 250 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=6480 $D=0
M2210 674 668 251 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=11110 $D=0
M2211 255 675 672 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=1850 $D=0
M2212 256 676 673 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=6480 $D=0
M2213 257 677 674 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=11110 $D=0
M2214 675 108 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=1850 $D=0
M2215 676 108 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=6480 $D=0
M2216 677 108 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=11110 $D=0
M2217 167 109 678 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=1850 $D=0
M2218 173 109 679 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=6480 $D=0
M2219 174 109 680 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=11110 $D=0
M2220 681 110 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=1850 $D=0
M2221 682 110 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=6480 $D=0
M2222 683 110 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=11110 $D=0
M2223 684 678 234 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=1850 $D=0
M2224 685 679 235 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=6480 $D=0
M2225 686 680 236 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=11110 $D=0
M2226 167 684 1044 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=1850 $D=0
M2227 173 685 1045 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=6480 $D=0
M2228 174 686 1046 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=11110 $D=0
M2229 687 1044 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=1850 $D=0
M2230 688 1045 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=6480 $D=0
M2231 689 1046 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=11110 $D=0
M2232 684 109 687 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=1850 $D=0
M2233 685 109 688 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=6480 $D=0
M2234 686 109 689 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=11110 $D=0
M2235 687 681 249 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=1850 $D=0
M2236 688 682 250 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=6480 $D=0
M2237 689 683 251 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=11110 $D=0
M2238 255 690 687 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=1850 $D=0
M2239 256 691 688 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=6480 $D=0
M2240 257 692 689 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=11110 $D=0
M2241 690 111 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=1850 $D=0
M2242 691 111 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=6480 $D=0
M2243 692 111 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=11110 $D=0
M2244 167 112 693 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=1850 $D=0
M2245 173 112 694 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=6480 $D=0
M2246 174 112 695 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=11110 $D=0
M2247 696 113 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=1850 $D=0
M2248 697 113 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=6480 $D=0
M2249 698 113 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=11110 $D=0
M2250 699 693 234 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=1850 $D=0
M2251 700 694 235 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=6480 $D=0
M2252 701 695 236 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=11110 $D=0
M2253 167 699 1047 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=1850 $D=0
M2254 173 700 1048 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=6480 $D=0
M2255 174 701 1049 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=11110 $D=0
M2256 702 1047 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=1850 $D=0
M2257 703 1048 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=6480 $D=0
M2258 704 1049 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=11110 $D=0
M2259 699 112 702 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=1850 $D=0
M2260 700 112 703 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=6480 $D=0
M2261 701 112 704 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=11110 $D=0
M2262 702 696 249 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=1850 $D=0
M2263 703 697 250 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=6480 $D=0
M2264 704 698 251 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=11110 $D=0
M2265 255 705 702 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=1850 $D=0
M2266 256 706 703 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=6480 $D=0
M2267 257 707 704 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=11110 $D=0
M2268 705 114 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=1850 $D=0
M2269 706 114 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=6480 $D=0
M2270 707 114 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=11110 $D=0
M2271 167 115 708 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=1850 $D=0
M2272 173 115 709 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=6480 $D=0
M2273 174 115 710 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=11110 $D=0
M2274 711 116 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=1850 $D=0
M2275 712 116 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=6480 $D=0
M2276 713 116 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=11110 $D=0
M2277 7 711 249 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=1850 $D=0
M2278 8 712 250 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=6480 $D=0
M2279 9 713 251 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=11110 $D=0
M2280 255 708 7 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=1850 $D=0
M2281 256 709 8 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=6480 $D=0
M2282 257 710 9 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=11110 $D=0
M2283 167 717 714 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=1850 $D=0
M2284 173 718 715 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=6480 $D=0
M2285 174 719 716 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=11110 $D=0
M2286 717 117 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=1850 $D=0
M2287 718 117 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=6480 $D=0
M2288 719 117 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=11110 $D=0
M2289 1050 249 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=1850 $D=0
M2290 1051 250 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=6480 $D=0
M2291 1052 251 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=11110 $D=0
M2292 720 717 1050 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=1850 $D=0
M2293 721 718 1051 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=6480 $D=0
M2294 722 719 1052 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=11110 $D=0
M2295 167 720 118 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=1850 $D=0
M2296 173 721 723 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=6480 $D=0
M2297 174 722 724 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=11110 $D=0
M2298 1053 118 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=1850 $D=0
M2299 1054 723 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=6480 $D=0
M2300 1055 724 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=11110 $D=0
M2301 720 714 1053 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=1850 $D=0
M2302 721 715 1054 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=6480 $D=0
M2303 722 716 1055 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=11110 $D=0
M2304 167 728 725 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=1850 $D=0
M2305 173 729 726 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=6480 $D=0
M2306 174 730 727 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=11110 $D=0
M2307 728 117 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=1850 $D=0
M2308 729 117 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=6480 $D=0
M2309 730 117 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=11110 $D=0
M2310 1056 255 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=1850 $D=0
M2311 1057 256 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=6480 $D=0
M2312 1058 257 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=11110 $D=0
M2313 731 728 1056 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=1850 $D=0
M2314 732 729 1057 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=6480 $D=0
M2315 733 730 1058 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=11110 $D=0
M2316 167 731 119 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=1850 $D=0
M2317 173 732 120 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=6480 $D=0
M2318 174 733 121 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=11110 $D=0
M2319 1059 119 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=1850 $D=0
M2320 1060 120 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=6480 $D=0
M2321 1061 121 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=11110 $D=0
M2322 731 725 1059 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=1850 $D=0
M2323 732 726 1060 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=6480 $D=0
M2324 733 727 1061 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=11110 $D=0
M2325 734 122 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=1850 $D=0
M2326 735 122 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=6480 $D=0
M2327 736 122 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=11110 $D=0
M2328 737 122 118 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=1850 $D=0
M2329 738 122 723 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=6480 $D=0
M2330 739 122 724 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=11110 $D=0
M2331 123 734 737 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=1850 $D=0
M2332 124 735 738 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=6480 $D=0
M2333 125 736 739 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=11110 $D=0
M2334 740 126 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=1850 $D=0
M2335 741 126 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=6480 $D=0
M2336 742 126 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=11110 $D=0
M2337 743 126 119 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=1850 $D=0
M2338 744 126 120 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=6480 $D=0
M2339 745 126 121 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=11110 $D=0
M2340 1062 740 743 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=1850 $D=0
M2341 1063 741 744 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=6480 $D=0
M2342 1064 742 745 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=11110 $D=0
M2343 167 119 1062 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=1850 $D=0
M2344 173 120 1063 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=6480 $D=0
M2345 174 121 1064 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=11110 $D=0
M2346 746 127 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=1850 $D=0
M2347 747 127 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=6480 $D=0
M2348 748 127 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=11110 $D=0
M2349 749 127 743 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=1850 $D=0
M2350 750 127 744 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=6480 $D=0
M2351 751 127 745 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=11110 $D=0
M2352 14 746 749 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=1850 $D=0
M2353 15 747 750 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=6480 $D=0
M2354 16 748 751 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=11110 $D=0
M2355 755 752 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=1850 $D=0
M2356 756 753 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=6480 $D=0
M2357 757 754 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=11110 $D=0
M2358 167 761 758 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=1850 $D=0
M2359 173 762 759 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=6480 $D=0
M2360 174 763 760 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=11110 $D=0
M2361 764 737 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=1850 $D=0
M2362 765 738 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=6480 $D=0
M2363 766 739 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=11110 $D=0
M2364 761 737 752 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=1850 $D=0
M2365 762 738 753 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=6480 $D=0
M2366 763 739 754 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=11110 $D=0
M2367 755 764 761 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=1850 $D=0
M2368 756 765 762 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=6480 $D=0
M2369 757 766 763 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=11110 $D=0
M2370 767 758 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=1850 $D=0
M2371 768 759 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=6480 $D=0
M2372 769 760 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=11110 $D=0
M2373 770 758 749 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=1850 $D=0
M2374 771 759 750 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=6480 $D=0
M2375 772 760 751 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=11110 $D=0
M2376 737 767 770 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=1850 $D=0
M2377 738 768 771 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=6480 $D=0
M2378 739 769 772 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=11110 $D=0
M2379 773 770 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=1850 $D=0
M2380 774 771 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=6480 $D=0
M2381 775 772 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=11110 $D=0
M2382 776 758 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=1850 $D=0
M2383 777 759 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=6480 $D=0
M2384 778 760 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=11110 $D=0
M2385 779 758 773 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=1850 $D=0
M2386 780 759 774 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=6480 $D=0
M2387 781 760 775 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=11110 $D=0
M2388 749 776 779 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=1850 $D=0
M2389 750 777 780 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=6480 $D=0
M2390 751 778 781 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=11110 $D=0
M2391 1095 737 167 167 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=1490 $D=0
M2392 1096 738 173 173 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=6120 $D=0
M2393 1097 739 174 174 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=10750 $D=0
M2394 782 749 1095 167 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=1490 $D=0
M2395 783 750 1096 173 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=6120 $D=0
M2396 784 751 1097 174 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=10750 $D=0
M2397 785 779 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=1850 $D=0
M2398 786 780 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=6480 $D=0
M2399 787 781 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=11110 $D=0
M2400 788 737 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=1850 $D=0
M2401 789 738 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=6480 $D=0
M2402 790 739 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=11110 $D=0
M2403 167 749 788 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=1850 $D=0
M2404 173 750 789 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=6480 $D=0
M2405 174 751 790 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=11110 $D=0
M2406 791 737 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=1850 $D=0
M2407 792 738 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=6480 $D=0
M2408 793 739 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=11110 $D=0
M2409 167 749 791 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=1850 $D=0
M2410 173 750 792 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=6480 $D=0
M2411 174 751 793 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=11110 $D=0
M2412 1098 737 167 167 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=1670 $D=0
M2413 1099 738 173 173 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=6300 $D=0
M2414 1100 739 174 174 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=10930 $D=0
M2415 797 749 1098 167 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=1670 $D=0
M2416 798 750 1099 173 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=6300 $D=0
M2417 799 751 1100 174 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=10930 $D=0
M2418 167 791 797 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=1850 $D=0
M2419 173 792 798 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=6480 $D=0
M2420 174 793 799 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=11110 $D=0
M2421 800 131 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=1850 $D=0
M2422 801 131 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=6480 $D=0
M2423 802 131 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=11110 $D=0
M2424 803 131 782 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=1850 $D=0
M2425 804 131 783 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=6480 $D=0
M2426 805 131 784 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=11110 $D=0
M2427 788 800 803 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=1850 $D=0
M2428 789 801 804 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=6480 $D=0
M2429 790 802 805 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=11110 $D=0
M2430 806 131 785 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=1850 $D=0
M2431 807 131 786 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=6480 $D=0
M2432 808 131 787 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=11110 $D=0
M2433 797 800 806 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=1850 $D=0
M2434 798 801 807 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=6480 $D=0
M2435 799 802 808 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=11110 $D=0
M2436 809 132 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=1850 $D=0
M2437 810 132 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=6480 $D=0
M2438 811 132 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=11110 $D=0
M2439 812 132 806 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=1850 $D=0
M2440 813 132 807 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=6480 $D=0
M2441 814 132 808 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=11110 $D=0
M2442 803 809 812 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=1850 $D=0
M2443 804 810 813 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=6480 $D=0
M2444 805 811 814 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=11110 $D=0
M2445 17 812 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=1850 $D=0
M2446 18 813 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=6480 $D=0
M2447 19 814 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=11110 $D=0
M2448 815 133 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=1850 $D=0
M2449 816 133 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=6480 $D=0
M2450 817 133 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=11110 $D=0
M2451 818 133 134 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=1850 $D=0
M2452 819 133 135 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=6480 $D=0
M2453 820 133 136 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=11110 $D=0
M2454 137 815 818 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=1850 $D=0
M2455 138 816 819 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=6480 $D=0
M2456 134 817 820 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=11110 $D=0
M2457 821 133 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=1850 $D=0
M2458 822 133 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=6480 $D=0
M2459 823 133 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=11110 $D=0
M2460 830 133 139 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=1850 $D=0
M2461 831 133 140 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=6480 $D=0
M2462 832 133 141 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=11110 $D=0
M2463 137 821 830 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=1850 $D=0
M2464 137 822 831 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=6480 $D=0
M2465 142 823 832 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=11110 $D=0
M2466 833 133 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=1850 $D=0
M2467 834 133 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=6480 $D=0
M2468 835 133 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=11110 $D=0
M2469 836 133 130 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=1850 $D=0
M2470 837 133 129 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=6480 $D=0
M2471 838 133 128 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=11110 $D=0
M2472 137 833 836 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=1850 $D=0
M2473 137 834 837 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=6480 $D=0
M2474 137 835 838 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=11110 $D=0
M2475 839 133 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=1850 $D=0
M2476 840 133 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=6480 $D=0
M2477 841 133 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=11110 $D=0
M2478 842 133 143 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=1850 $D=0
M2479 843 133 144 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=6480 $D=0
M2480 844 133 145 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=11110 $D=0
M2481 137 839 842 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=1850 $D=0
M2482 137 840 843 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=6480 $D=0
M2483 137 841 844 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=11110 $D=0
M2484 845 133 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=1850 $D=0
M2485 846 133 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=6480 $D=0
M2486 847 133 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=11110 $D=0
M2487 848 133 146 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=1850 $D=0
M2488 849 133 147 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=6480 $D=0
M2489 850 133 148 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=11110 $D=0
M2490 137 845 848 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=1850 $D=0
M2491 137 846 849 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=6480 $D=0
M2492 137 847 850 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=11110 $D=0
M2493 167 737 1080 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=1850 $D=0
M2494 173 738 1081 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=6480 $D=0
M2495 174 739 1082 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=11110 $D=0
M2496 138 1080 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=1850 $D=0
M2497 134 1081 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=6480 $D=0
M2498 135 1082 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=11110 $D=0
M2499 851 149 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=1850 $D=0
M2500 852 149 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=6480 $D=0
M2501 853 149 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=11110 $D=0
M2502 150 149 138 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=1850 $D=0
M2503 151 149 134 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=6480 $D=0
M2504 139 149 135 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=11110 $D=0
M2505 818 851 150 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=1850 $D=0
M2506 819 852 151 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=6480 $D=0
M2507 820 853 139 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=11110 $D=0
M2508 854 152 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=1850 $D=0
M2509 855 152 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=6480 $D=0
M2510 856 152 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=11110 $D=0
M2511 153 152 150 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=1850 $D=0
M2512 154 152 151 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=6480 $D=0
M2513 155 152 139 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=11110 $D=0
M2514 830 854 153 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=1850 $D=0
M2515 831 855 154 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=6480 $D=0
M2516 832 856 155 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=11110 $D=0
M2517 857 156 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=1850 $D=0
M2518 858 156 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=6480 $D=0
M2519 859 156 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=11110 $D=0
M2520 157 156 153 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=1850 $D=0
M2521 158 156 154 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=6480 $D=0
M2522 159 156 155 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=11110 $D=0
M2523 836 857 157 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=1850 $D=0
M2524 837 858 158 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=6480 $D=0
M2525 838 859 159 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=11110 $D=0
M2526 860 160 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=1850 $D=0
M2527 861 160 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=6480 $D=0
M2528 862 160 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=11110 $D=0
M2529 161 160 157 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=1850 $D=0
M2530 162 160 158 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=6480 $D=0
M2531 163 160 159 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=11110 $D=0
M2532 842 860 161 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=1850 $D=0
M2533 843 861 162 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=6480 $D=0
M2534 844 862 163 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=11110 $D=0
M2535 863 164 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=1850 $D=0
M2536 864 164 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=6480 $D=0
M2537 865 164 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=11110 $D=0
M2538 213 164 161 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=1850 $D=0
M2539 214 164 162 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=6480 $D=0
M2540 215 164 163 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=11110 $D=0
M2541 848 863 213 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=1850 $D=0
M2542 849 864 214 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=6480 $D=0
M2543 850 865 215 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=11110 $D=0
M2544 866 165 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=1850 $D=0
M2545 867 165 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=6480 $D=0
M2546 868 165 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=11110 $D=0
M2547 166 165 119 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=1850 $D=0
M2548 869 165 120 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=6480 $D=0
M2549 870 165 121 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=11110 $D=0
M2550 14 866 166 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=1850 $D=0
M2551 15 867 869 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=6480 $D=0
M2552 16 868 870 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=11110 $D=0
M2553 871 118 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=1850 $D=0
M2554 872 723 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=6480 $D=0
M2555 873 724 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=11110 $D=0
M2556 167 166 871 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=1850 $D=0
M2557 173 869 872 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=6480 $D=0
M2558 174 870 873 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=11110 $D=0
M2559 1101 118 167 167 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=1670 $D=0
M2560 1102 723 173 173 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=6300 $D=0
M2561 1103 724 174 174 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=10930 $D=0
M2562 877 166 1101 167 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=1670 $D=0
M2563 878 869 1102 173 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=6300 $D=0
M2564 879 870 1103 174 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=10930 $D=0
M2565 167 871 877 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=1850 $D=0
M2566 173 872 878 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=6480 $D=0
M2567 174 873 879 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=11110 $D=0
M2568 1083 167 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=1850 $D=0
M2569 1084 880 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=6480 $D=0
M2570 1085 881 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=11110 $D=0
M2571 167 877 1083 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=1850 $D=0
M2572 173 878 1084 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=6480 $D=0
M2573 174 879 1085 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=11110 $D=0
M2574 880 1083 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=1850 $D=0
M2575 881 1084 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=6480 $D=0
M2576 168 1085 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=11110 $D=0
M2577 1104 118 167 167 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=1490 $D=0
M2578 1105 723 173 173 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=6120 $D=0
M2579 1106 724 174 174 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=10750 $D=0
M2580 882 885 1104 167 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=1490 $D=0
M2581 883 886 1105 173 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=6120 $D=0
M2582 884 887 1106 174 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=10750 $D=0
M2583 885 166 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=1850 $D=0
M2584 886 869 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=6480 $D=0
M2585 887 870 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=11110 $D=0
M2586 888 882 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=1850 $D=0
M2587 889 883 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=6480 $D=0
M2588 890 884 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=11110 $D=0
M2589 167 167 888 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=1850 $D=0
M2590 173 880 889 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=6480 $D=0
M2591 174 881 890 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=11110 $D=0
M2592 893 7 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=1850 $D=0
M2593 894 891 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=6480 $D=0
M2594 895 892 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=11110 $D=0
M2595 891 888 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=1850 $D=0
M2596 892 889 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=6480 $D=0
M2597 169 890 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=11110 $D=0
M2598 167 893 891 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=1850 $D=0
M2599 173 894 892 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=6480 $D=0
M2600 174 895 169 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=11110 $D=0
M2601 898 896 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=1850 $D=0
M2602 899 897 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=6480 $D=0
M2603 900 170 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=11110 $D=0
M2604 167 904 901 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=1850 $D=0
M2605 173 905 902 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=6480 $D=0
M2606 174 906 903 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=11110 $D=0
M2607 907 123 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=1850 $D=0
M2608 908 124 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=6480 $D=0
M2609 909 125 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=11110 $D=0
M2610 904 123 896 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=1850 $D=0
M2611 905 124 897 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=6480 $D=0
M2612 906 125 170 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=11110 $D=0
M2613 898 907 904 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=1850 $D=0
M2614 899 908 905 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=6480 $D=0
M2615 900 909 906 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=11110 $D=0
M2616 910 901 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=1850 $D=0
M2617 911 902 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=6480 $D=0
M2618 912 903 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=11110 $D=0
M2619 913 901 7 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=1850 $D=0
M2620 896 902 8 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=6480 $D=0
M2621 897 903 9 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=11110 $D=0
M2622 123 910 913 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=1850 $D=0
M2623 124 911 896 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=6480 $D=0
M2624 125 912 897 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=11110 $D=0
M2625 914 913 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=1850 $D=0
M2626 915 896 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=6480 $D=0
M2627 916 897 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=11110 $D=0
M2628 917 901 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=1850 $D=0
M2629 918 902 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=6480 $D=0
M2630 919 903 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=11110 $D=0
M2631 216 901 914 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=1850 $D=0
M2632 217 902 915 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=6480 $D=0
M2633 218 903 916 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=11110 $D=0
M2634 7 917 216 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=1850 $D=0
M2635 8 918 217 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=6480 $D=0
M2636 9 919 218 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=11110 $D=0
M2637 920 171 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=1850 $D=0
M2638 921 171 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=6480 $D=0
M2639 922 171 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=11110 $D=0
M2640 923 171 216 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=1850 $D=0
M2641 924 171 217 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=6480 $D=0
M2642 925 171 218 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=11110 $D=0
M2643 17 920 923 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=1850 $D=0
M2644 18 921 924 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=6480 $D=0
M2645 19 922 925 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=11110 $D=0
M2646 926 172 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=1850 $D=0
M2647 927 172 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=6480 $D=0
M2648 928 172 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=11110 $D=0
M2649 929 172 923 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=1850 $D=0
M2650 172 172 924 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=6480 $D=0
M2651 172 172 925 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=11110 $D=0
M2652 7 926 929 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=1850 $D=0
M2653 173 927 172 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=6480 $D=0
M2654 174 928 172 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=11110 $D=0
M2655 930 117 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=1850 $D=0
M2656 931 117 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=6480 $D=0
M2657 932 117 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=11110 $D=0
M2658 167 930 933 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=1850 $D=0
M2659 173 931 934 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=6480 $D=0
M2660 174 932 935 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=11110 $D=0
M2661 936 117 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=1850 $D=0
M2662 937 117 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=6480 $D=0
M2663 938 117 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=11110 $D=0
M2664 939 933 929 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=1850 $D=0
M2665 940 934 172 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=6480 $D=0
M2666 941 935 172 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=11110 $D=0
M2667 167 939 1086 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=1850 $D=0
M2668 173 940 1087 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=6480 $D=0
M2669 174 941 1088 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=11110 $D=0
M2670 942 1086 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=1850 $D=0
M2671 943 1087 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=6480 $D=0
M2672 944 1088 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=11110 $D=0
M2673 939 930 942 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=1850 $D=0
M2674 940 931 943 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=6480 $D=0
M2675 941 932 944 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=11110 $D=0
M2676 945 936 942 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=1850 $D=0
M2677 946 937 943 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=6480 $D=0
M2678 947 938 944 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=11110 $D=0
M2679 167 951 948 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=1850 $D=0
M2680 173 952 949 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=6480 $D=0
M2681 174 953 950 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=11110 $D=0
M2682 951 117 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=1850 $D=0
M2683 952 117 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=6480 $D=0
M2684 953 117 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=11110 $D=0
M2685 1089 945 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=1850 $D=0
M2686 1090 946 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=6480 $D=0
M2687 1091 947 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=11110 $D=0
M2688 954 951 1089 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=1850 $D=0
M2689 955 952 1090 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=6480 $D=0
M2690 956 953 1091 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=11110 $D=0
M2691 167 954 123 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=1850 $D=0
M2692 173 955 124 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=6480 $D=0
M2693 174 956 125 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=11110 $D=0
M2694 1092 123 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=1850 $D=0
M2695 1093 124 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=6480 $D=0
M2696 1094 125 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=11110 $D=0
M2697 954 948 1092 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=1850 $D=0
M2698 955 949 1093 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=6480 $D=0
M2699 956 950 1094 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=11110 $D=0
.ENDS
***************************************
.SUBCKT datapath 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 vss! vdd!
+ 61 62 63 64 shift_out<114> mem_mux_sel<0> dmem_rdata<2> dmem_rdata<1> dmem_rdata<0> mem_mux_sel<1> mem_mux_sel<2> rd_mux_sel<0> cmp_out imm<2> imm<1> imm<0> rd_mux_sel<1> rd_mux_sel<2> rd_sel<31> rs1_sel<31>
+ rs2_sel<31> rd_sel<30> rs1_sel<30> rs2_sel<30> rd_sel<29> rs1_sel<29> rs2_sel<29> rd_sel<28> rs1_sel<28> rs2_sel<28> rd_sel<27> rs1_sel<27> rs2_sel<27> rd_sel<26> rs1_sel<26> rs2_sel<26> rd_sel<25> rs1_sel<25> rs2_sel<25> rd_sel<24>
+ rs1_sel<24> rs2_sel<24> rd_sel<23> rs1_sel<23> rs2_sel<23> rd_sel<22> rs1_sel<22> rs2_sel<22> rd_sel<21> rs1_sel<21> rs2_sel<21> rd_sel<20> rs1_sel<20> rs2_sel<20> rd_sel<19> rs1_sel<19> rs2_sel<19> rd_sel<18> rs1_sel<18> rs2_sel<18>
+ rd_sel<17> rs1_sel<17> rs2_sel<17> rd_sel<16> rs1_sel<16> rs2_sel<16> rd_sel<15> rs1_sel<15> rs2_sel<15> rd_sel<14> rs1_sel<14> rs2_sel<14> rd_sel<13> rs1_sel<13> rs2_sel<13> rd_sel<12> rs1_sel<12> rs2_sel<12> rd_sel<11> rs1_sel<11>
+ rs2_sel<11> rd_sel<10> rs1_sel<10> rs2_sel<10> rd_sel<9> rs1_sel<9> rs2_sel<9> rd_sel<8> rs1_sel<8> rs2_sel<8> rd_sel<7> rs1_sel<7> rs2_sel<7> rd_sel<6> rs1_sel<6> rs2_sel<6> rd_sel<5> rs1_sel<5> rs2_sel<5> rd_sel<4>
+ rs1_sel<4> rs2_sel<4> rd_sel<3> rs1_sel<3> rs2_sel<3> rd_sel<2> rs1_sel<2> rs2_sel<2> rd_sel<1> rs1_sel<1> rs2_sel<1> rs2_sel<0> rs1_sel<0> clk dmem_wdata<2> dmem_wdata<1> dmem_wdata<0> alu_mux_1_sel alu_inv_rs2 alu_mux_2_sel
+ alu_cin shift_out<2> shift_out<7> shift_out<12> alu_op<0> alu_op<1> shift_out<16> dmem_addr<2> dmem_addr<1> dmem_addr<0> shift_dir shift_amount<2> shift_amount<1> shift_out<0> shift_out<15> shift_out<6> shift_out<1> shift_out<21> shift_out<11> shift_out<32>
+ shift_out<27> shift_out<22> shift_out<53> shift_out<48> shift_out<43> shift_out<94> shift_out<89> shift_amount<3> 216 217 218 shift_amount<4> 220 221 222 cmp_mux_sel cmp_eq cmp_lt pc_mux_sel rst
+ imem_addr<2> imem_addr<1> imem_addr<0> dmem_rdata<4> dmem_rdata<3> imm<4> imm<3> dmem_wdata<4> dmem_wdata<3> shift_out<17> 242 shift_out<26> dmem_addr<3> dmem_addr<4> shift_out<25> shift_out<31> shift_out<37> shift_out<63> shift_out<58> shift_out<104>
+ shift_out<99> 253 254 255 256 imem_addr<4> imem_addr<3> dmem_rdata<6> dmem_rdata<5> imm<6> imm<5> dmem_wdata<6> dmem_wdata<5> shift_out<36> dmem_addr<6> dmem_addr<5> shift_out<30> shift_out<35> shift_out<41> shift_out<52>
+ shift_out<47> shift_out<73> shift_out<68> shift_out<109> 280 281 282 283 imem_addr<6> imem_addr<5> dmem_rdata<8> dmem_rdata<7> imm<8> imm<7> dmem_wdata<8> dmem_wdata<7> shift_out<46> dmem_addr<8> dmem_addr<7> shift_out<40>
+ shift_out<45> shift_out<51> 302 303 shift_out<3> 305 306 shift_out<124> shift_out<119> 309 310 311 312 imem_addr<8> imem_addr<7> dmem_rdata<10> dmem_rdata<9> imm<10> imm<9> dmem_wdata<10>
+ dmem_wdata<9> shift_out<56> dmem_addr<9> dmem_addr<10> shift_out<50> shift_out<55> shift_out<61> 331 332 333 334 shift_out<13> shift_out<8> 337 338 shift_out<134> shift_out<129> 341 342 imem_addr<10>
+ imem_addr<9> dmem_rdata<12> dmem_rdata<11> imm<12> imm<11> dmem_wdata<12> dmem_wdata<11> shift_out<62> shift_out<66> dmem_addr<11> dmem_addr<12> shift_out<60> shift_out<65> shift_out<71> shift_out<42> 363 364 365 shift_out<23> shift_out<18>
+ 368 shift_out<98> shift_out<144> shift_out<139> 372 373 374 imem_addr<12> imem_addr<11> dmem_rdata<14> dmem_rdata<13> imm<14> imm<13> dmem_wdata<14> dmem_wdata<13> shift_out<67> shift_out<72> shift_out<76> dmem_addr<14> dmem_addr<13>
+ shift_out<70> shift_out<75> shift_out<81> 395 396 397 398 shift_out<33> shift_out<28> 401 402 shift_out<154> shift_out<149> 405 406 imem_addr<14> imem_addr<13> dmem_rdata<16> dmem_rdata<15> imm<16>
+ imm<15> dmem_wdata<16> dmem_wdata<15> shift_out<82> shift_out<77> shift_out<86> dmem_addr<16> dmem_addr<15> shift_out<80> shift_out<91> shift_out<57> 427 428 429 shift_out<38> shift_out<123> 432 shift_out<4> shift_msb shift_out<159>
+ shift_out<85> 437 438 shift_out<84> 440 imem_addr<16> imem_addr<15> dmem_rdata<20> dmem_rdata<19> dmem_rdata<18> dmem_rdata<17> imm<20> imm<19> imm<18> imm<17> dmem_wdata<20> dmem_wdata<19> dmem_wdata<18> dmem_wdata<17> shift_out<87>
+ shift_out<92> shift_out<97> shift_out<96> shift_out<106> dmem_addr<17> dmem_addr<20> dmem_addr<19> dmem_addr<18> shift_out<95> shift_out<90> shift_out<105> shift_out<100> shift_out<111> shift_out<101> 474 475 476 477 478 479
+ 480 481 shift_out<143> shift_out<138> shift_out<133> shift_out<128> shift_out<24> shift_out<19> shift_out<14> shift_out<9> shift_out<102> 491 492 493 494 495 496 497 498 imem_addr<20>
+ imem_addr<19> imem_addr<18> imem_addr<17> dmem_rdata<22> dmem_rdata<21> imm<22> imm<21> dmem_wdata<22> dmem_wdata<21> shift_out<107> shift_out<116> dmem_addr<22> dmem_addr<21> shift_out<115> shift_out<110> shift_out<121> 520 521 522 523
+ shift_out<153> shift_out<148> shift_out<34> shift_out<29> shift_out<112> 529 530 531 532 imem_addr<22> imem_addr<21> dmem_rdata<24> dmem_rdata<23> imm<24> imm<23> dmem_wdata<24> dmem_wdata<23> shift_out<117> shift_out<126> dmem_addr<24>
+ dmem_addr<23> shift_out<125> shift_out<120> shift_out<131> shift_out<142> 552 shift_out<83> shift_out<78> shift_out<158> shift_out<44> shift_out<39> shift_out<122> 559 560 561 562 imem_addr<24> imem_addr<23> dmem_rdata<26> dmem_rdata<25>
+ imm<26> imm<25> dmem_wdata<26> dmem_wdata<25> shift_out<127> shift_out<136> dmem_addr<26> dmem_addr<25> shift_out<135> shift_out<130> shift_out<141> shift_out<152> shift_out<147> shift_out<93> shift_out<88> shift_out<54> shift_out<49> shift_out<132> 588 589
+ 590 591 imem_addr<26> imem_addr<25> dmem_rdata<28> dmem_rdata<27> imm<28> imm<27> dmem_wdata<28> dmem_wdata<27> shift_out<137> shift_out<146> dmem_addr<28> dmem_addr<27> shift_out<145> shift_out<140> shift_out<151> shift_out<157> shift_out<103> shift_out98>
+ shift_out<64> shift_out<59> 616 617 618 619 620 imem_addr<28> imem_addr<27> dmem_rdata<31> dmem_rdata<30> dmem_rdata<29> imm<31> imm<30> imm<29> dmem_wdata<31> dmem_wdata<30> dmem_wdata<29> dmem_addr<31> dmem_addr<30>
+ dmem_addr<29> shift_out<150> shift_out<155> shift_out<156> shift_out<118> shift_out<113> shift_out<108> shift_out<79> shift_out<74> shift_out<69> 646 647 648 649 650 651 652 653 654 655
+ cmp_a_31 cmp_b_31 imem_addr<31> imem_addr<30> imem_addr<29>
** N=660 EP=605 IP=2451 FDC=28800
X0 mem_mux_sel<0> dmem_rdata<2> dmem_rdata<1> dmem_rdata<0> mem_mux_sel<1> mem_mux_sel<2> rd_mux_sel<0> 1 3 cmp_out imm<2> imm<1> imm<0> dmem_addr<2> dmem_addr<1> dmem_addr<0> rd_mux_sel<1> rd_mux_sel<2> rd_sel<31> rs1_sel<31>
+ rs2_sel<31> rd_sel<30> rs1_sel<30> rs2_sel<30> rd_sel<29> rs1_sel<29> rs2_sel<29> rd_sel<28> rs1_sel<28> rs2_sel<28> rd_sel<27> rs1_sel<27> rs2_sel<27> rd_sel<26> rs1_sel<26> rs2_sel<26> rd_sel<25> rs1_sel<25> rs2_sel<25> rd_sel<24>
+ rs1_sel<24> rs2_sel<24> rd_sel<23> rs1_sel<23> rs2_sel<23> rd_sel<22> rs1_sel<22> rs2_sel<22> rd_sel<21> rs1_sel<21> rs2_sel<21> rd_sel<20> rs1_sel<20> rs2_sel<20> rd_sel<19> rs1_sel<19> rs2_sel<19> rd_sel<18> rs1_sel<18> rs2_sel<18>
+ rd_sel<17> rs1_sel<17> rs2_sel<17> rd_sel<16> rs1_sel<16> rs2_sel<16> rd_sel<15> rs1_sel<15> rs2_sel<15> rd_sel<14> rs1_sel<14> rs2_sel<14> rd_sel<13> rs1_sel<13> rs2_sel<13> rd_sel<12> rs1_sel<12> rs2_sel<12> rd_sel<11> rs1_sel<11>
+ rs2_sel<11> rd_sel<10> rs1_sel<10> rs2_sel<10> rd_sel<9> rs1_sel<9> rs2_sel<9> rd_sel<8> rs1_sel<8> rs2_sel<8> rd_sel<7> rs1_sel<7> rs2_sel<7> rd_sel<6> rs1_sel<6> rs2_sel<6> rd_sel<5> rs1_sel<5> rs2_sel<5> rd_sel<4>
+ rs1_sel<4> rs2_sel<4> rd_sel<3> rs1_sel<3> rs2_sel<3> rd_sel<2> rs1_sel<2> rs2_sel<2> rd_sel<1> rs1_sel<1> rs2_sel<1> rs2_sel<0> rs1_sel<0> clk dmem_wdata<2> dmem_wdata<1> dmem_wdata<0> alu_mux_1_sel imem_addr<2> imem_addr<1>
+ imem_addr<0> alu_inv_rs2 alu_mux_2_sel shift_amount<2> shift_amount<1> 214 alu_cin 186 shift_out<2> shift_out<7> shift_out<12> alu_op<0> alu_op<1> shift_dir shift_out<0> 5 shift_out<15> shift_out<1> shift_out<21> shift_out<16>
+ shift_out<11> shift_out<32> shift_out<27> shift_out<22> shift_out<53> shift_out<48> shift_out<43> shift_out<94> shift_out<89> shift_out<6> 216 217 218 shift_amount<3> 220 221 222 shift_amount<4> cmp_mux_sel cmp_eq
+ 226 cmp_lt 2 228 pc_mux_sel rst 4 6
+ ICV_24 $T=0 0 0 0 $X=0 $Y=132400
X1 mem_mux_sel<0> dmem_rdata<4> dmem_rdata<3> mem_mux_sel<1> mem_mux_sel<2> rd_mux_sel<0> 7 9 imm<4> imm<3> dmem_addr<4> dmem_addr<3> rd_mux_sel<1> rd_mux_sel<2> rd_sel<31> rs1_sel<31> rs2_sel<31> rd_sel<30> rs1_sel<30> rs2_sel<30>
+ rd_sel<29> rs1_sel<29> rs2_sel<29> rd_sel<28> rs1_sel<28> rs2_sel<28> rd_sel<27> rs1_sel<27> rs2_sel<27> rd_sel<26> rs1_sel<26> rs2_sel<26> rd_sel<25> rs1_sel<25> rs2_sel<25> rd_sel<24> rs1_sel<24> rs2_sel<24> rd_sel<23> rs1_sel<23>
+ rs2_sel<23> rd_sel<22> rs1_sel<22> rs2_sel<22> rd_sel<21> rs1_sel<21> rs2_sel<21> rd_sel<20> rs1_sel<20> rs2_sel<20> rd_sel<19> rs1_sel<19> rs2_sel<19> rd_sel<18> rs1_sel<18> rs2_sel<18> rd_sel<17> rs1_sel<17> rs2_sel<17> rd_sel<16>
+ rs1_sel<16> rs2_sel<16> rd_sel<15> rs1_sel<15> rs2_sel<15> rd_sel<14> rs1_sel<14> rs2_sel<14> rd_sel<13> rs1_sel<13> rs2_sel<13> rd_sel<12> rs1_sel<12> rs2_sel<12> rd_sel<11> rs1_sel<11> rs2_sel<11> rd_sel<10> rs1_sel<10> rs2_sel<10>
+ rd_sel<9> rs1_sel<9> rs2_sel<9> rd_sel<8> rs1_sel<8> rs2_sel<8> rd_sel<7> rs1_sel<7> rs2_sel<7> rd_sel<6> rs1_sel<6> rs2_sel<6> rd_sel<5> rs1_sel<5> rs2_sel<5> rd_sel<4> rs1_sel<4> rs2_sel<4> rd_sel<3> rs1_sel<3>
+ rs2_sel<3> rd_sel<2> rs1_sel<2> rs2_sel<2> rd_sel<1> rs1_sel<1> rs2_sel<1> rs2_sel<0> rs1_sel<0> clk dmem_wdata<4> dmem_wdata<3> alu_mux_1_sel imem_addr<4> imem_addr<3> alu_inv_rs2 alu_mux_2_sel shift_amount<4> shift_amount<3> 186
+ shift_out<2> shift_out<17> alu_op<0> alu_op<1> 242 shift_dir shift_out<15> shift_amount<2> shift_out<25> shift_out<11> shift_out<26> shift_out<6> shift_out<31> shift_out<53> shift_out<37> shift_out<63> shift_out<58> shift_out<104> shift_out<99> 214
+ shift_out<21> shift_out<16> shift_amount<1> shift_out<22> 253 254 255 256 cmp_mux_sel 224 258 226 228 259 pc_mux_sel rst 8 10
+ ICV_25 $T=0 0 0 0 $X=0 $Y=123200
X2 mem_mux_sel<0> dmem_rdata<6> dmem_rdata<5> mem_mux_sel<1> mem_mux_sel<2> rd_mux_sel<0> 11 13 imm<6> imm<5> dmem_addr<6> dmem_addr<5> rd_mux_sel<1> rd_mux_sel<2> rd_sel<31> rs1_sel<31> rs2_sel<31> rd_sel<30> rs1_sel<30> rs2_sel<30>
+ rd_sel<29> rs1_sel<29> rs2_sel<29> rd_sel<28> rs1_sel<28> rs2_sel<28> rd_sel<27> rs1_sel<27> rs2_sel<27> rd_sel<26> rs1_sel<26> rs2_sel<26> rd_sel<25> rs1_sel<25> rs2_sel<25> rd_sel<24> rs1_sel<24> rs2_sel<24> rd_sel<23> rs1_sel<23>
+ rs2_sel<23> rd_sel<22> rs1_sel<22> rs2_sel<22> rd_sel<21> rs1_sel<21> rs2_sel<21> rd_sel<20> rs1_sel<20> rs2_sel<20> rd_sel<19> rs1_sel<19> rs2_sel<19> rd_sel<18> rs1_sel<18> rs2_sel<18> rd_sel<17> rs1_sel<17> rs2_sel<17> rd_sel<16>
+ rs1_sel<16> rs2_sel<16> rd_sel<15> rs1_sel<15> rs2_sel<15> rd_sel<14> rs1_sel<14> rs2_sel<14> rd_sel<13> rs1_sel<13> rs2_sel<13> rd_sel<12> rs1_sel<12> rs2_sel<12> rd_sel<11> rs1_sel<11> rs2_sel<11> rd_sel<10> rs1_sel<10> rs2_sel<10>
+ rd_sel<9> rs1_sel<9> rs2_sel<9> rd_sel<8> rs1_sel<8> rs2_sel<8> rd_sel<7> rs1_sel<7> rs2_sel<7> rd_sel<6> rs1_sel<6> rs2_sel<6> rd_sel<5> rs1_sel<5> rs2_sel<5> rd_sel<4> rs1_sel<4> rs2_sel<4> rd_sel<3> rs1_sel<3>
+ rs2_sel<3> rd_sel<2> rs1_sel<2> rs2_sel<2> rd_sel<1> rs1_sel<1> rs2_sel<1> rs2_sel<0> rs1_sel<0> clk dmem_wdata<6> dmem_wdata<5> alu_mux_1_sel imem_addr<6> imem_addr<5> alu_inv_rs2 alu_mux_2_sel 240 268 shift_out<12>
+ alu_op<0> alu_op<1> shift_dir shift_out<25> shift_amount<4> shift_out<35> shift_out<30> shift_out<21> shift_out<36> shift_out<16> shift_out<41> shift_out<7> shift_out<53> shift_out<52> shift_out<47> shift_out<73> shift_out<68> shift_out<114> shift_out<109> 214
+ shift_out<31> shift_out<26> shift_amount<1> shift_out<32> shift_out<27> shift_amount<2> 280 281 shift_amount<3> 282 283 cmp_mux_sel 257 285 258 259 286 pc_mux_sel rst 12
+ 14
+ ICV_26 $T=0 0 0 0 $X=0 $Y=114000
X3 mem_mux_sel<0> dmem_rdata<8> dmem_rdata<7> 15 mem_mux_sel<1> mem_mux_sel<2> rd_mux_sel<0> 17 imm<8> imm<7> dmem_addr<8> dmem_addr<7> rd_mux_sel<1> rd_mux_sel<2> rd_sel<31> rs1_sel<31> rs2_sel<31> rd_sel<30> rs1_sel<30> rs2_sel<30>
+ rd_sel<29> rs1_sel<29> rs2_sel<29> rd_sel<28> rs1_sel<28> rs2_sel<28> rd_sel<27> rs1_sel<27> rs2_sel<27> rd_sel<26> rs1_sel<26> rs2_sel<26> rd_sel<25> rs1_sel<25> rs2_sel<25> rd_sel<24> rs1_sel<24> rs2_sel<24> rd_sel<23> rs1_sel<23>
+ rs2_sel<23> rd_sel<22> rs1_sel<22> rs2_sel<22> rd_sel<21> rs1_sel<21> rs2_sel<21> rd_sel<20> rs1_sel<20> rs2_sel<20> rd_sel<19> rs1_sel<19> rs2_sel<19> rd_sel<18> rs1_sel<18> rs2_sel<18> rd_sel<17> rs1_sel<17> rs2_sel<17> rd_sel<16>
+ rs1_sel<16> rs2_sel<16> rd_sel<15> rs1_sel<15> rs2_sel<15> rd_sel<14> rs1_sel<14> rs2_sel<14> rd_sel<13> rs1_sel<13> rs2_sel<13> rd_sel<12> rs1_sel<12> rs2_sel<12> rd_sel<11> rs1_sel<11> rs2_sel<11> rd_sel<10> rs1_sel<10> rs2_sel<10>
+ rd_sel<9> rs1_sel<9> rs2_sel<9> rd_sel<8> rs1_sel<8> rs2_sel<8> rd_sel<7> rs1_sel<7> rs2_sel<7> rd_sel<6> rs1_sel<6> rs2_sel<6> rd_sel<5> rs1_sel<5> rs2_sel<5> rd_sel<4> rs1_sel<4> rs2_sel<4> rd_sel<3> rs1_sel<3>
+ rs2_sel<3> rd_sel<2> rs1_sel<2> rs2_sel<2> rd_sel<1> rs1_sel<1> rs2_sel<1> rs2_sel<0> rs1_sel<0> clk dmem_wdata<8> dmem_wdata<7> alu_mux_1_sel imem_addr<8> imem_addr<7> alu_inv_rs2 alu_mux_2_sel 268 alu_op<0> alu_op<1>
+ shift_dir shift_out<35> shift_out<30> shift_out<45> shift_out<40> 309 shift_out<31> shift_out<46> shift_out<26> shift_out<51> shift_out<22> shift_out<17> shift_out<53> 302 303 shift_out<3> 305 306 shift_out<124> shift_out<119>
+ 214 shift_out<43> shift_out<41> shift_out<36> shift_amount<1> shift_out<37> shift_amount<2> 310 shift_amount<3> 311 312 shift_amount<4> cmp_mux_sel 284 314 285 286 315 pc_mux_sel rst
+ 16 18
+ ICV_27 $T=0 0 0 0 $X=0 $Y=104600
X4 mem_mux_sel<0> dmem_rdata<10> dmem_rdata<9> dmem_rdata<7> 19 21 mem_mux_sel<1> mem_mux_sel<2> rd_mux_sel<0> imm<10> imm<9> dmem_addr<10> dmem_addr<9> rd_mux_sel<1> rd_mux_sel<2> rd_sel<31> rs1_sel<31> rs2_sel<31> rd_sel<30> rs1_sel<30>
+ rs2_sel<30> rd_sel<29> rs1_sel<29> rs2_sel<29> rd_sel<28> rs1_sel<28> rs2_sel<28> rd_sel<27> rs1_sel<27> rs2_sel<27> rd_sel<26> rs1_sel<26> rs2_sel<26> rd_sel<25> rs1_sel<25> rs2_sel<25> rd_sel<24> rs1_sel<24> rs2_sel<24> rd_sel<23>
+ rs1_sel<23> rs2_sel<23> rd_sel<22> rs1_sel<22> rs2_sel<22> rd_sel<21> rs1_sel<21> rs2_sel<21> rd_sel<20> rs1_sel<20> rs2_sel<20> rd_sel<19> rs1_sel<19> rs2_sel<19> rd_sel<18> rs1_sel<18> rs2_sel<18> rd_sel<17> rs1_sel<17> rs2_sel<17>
+ rd_sel<16> rs1_sel<16> rs2_sel<16> rd_sel<15> rs1_sel<15> rs2_sel<15> rd_sel<14> rs1_sel<14> rs2_sel<14> rd_sel<13> rs1_sel<13> rs2_sel<13> rd_sel<12> rs1_sel<12> rs2_sel<12> rd_sel<11> rs1_sel<11> rs2_sel<11> rd_sel<10> rs1_sel<10>
+ rs2_sel<10> rd_sel<9> rs1_sel<9> rs2_sel<9> rd_sel<8> rs1_sel<8> rs2_sel<8> rd_sel<7> rs1_sel<7> rs2_sel<7> rd_sel<6> rs1_sel<6> rs2_sel<6> rd_sel<5> rs1_sel<5> rs2_sel<5> rd_sel<4> rs1_sel<4> rs2_sel<4> rd_sel<3>
+ rs1_sel<3> rs2_sel<3> rd_sel<2> rs1_sel<2> rs2_sel<2> rd_sel<1> rs1_sel<1> rs2_sel<1> rs2_sel<0> rs1_sel<0> clk dmem_wdata<10> dmem_wdata<9> alu_mux_1_sel imem_addr<10> imem_addr<9> alu_inv_rs2 alu_mux_2_sel 295 324
+ alu_op<0> alu_op<1> shift_dir shift_out<45> shift_out<40> shift_out<55> shift_out<50> shift_out<41> shift_out<56> shift_out<36> shift_out<61> 331 332 shift_out<53> 333 334 shift_out<13> shift_out<8> 337 338
+ shift_out<134> shift_out<129> 214 shift_out<51> shift_out<46> shift_amount<1> shift_out<52> shift_out<47> shift_amount<2> shift_out<48> shift_amount<3> 341 342 shift_amount<4> cmp_mux_sel 313 344 314 315 345
+ pc_mux_sel rst 20 22
+ ICV_28 $T=0 0 0 0 $X=0 $Y=95400
X5 mem_mux_sel<0> dmem_rdata<12> dmem_rdata<11> dmem_rdata<7> 23 25 mem_mux_sel<1> mem_mux_sel<2> rd_mux_sel<0> imm<12> imm<11> dmem_addr<12> dmem_addr<11> rd_mux_sel<1> rd_mux_sel<2> rd_sel<31> rs1_sel<31> rs2_sel<31> rd_sel<30> rs1_sel<30>
+ rs2_sel<30> rd_sel<29> rs1_sel<29> rs2_sel<29> rd_sel<28> rs1_sel<28> rs2_sel<28> rd_sel<27> rs1_sel<27> rs2_sel<27> rd_sel<26> rs1_sel<26> rs2_sel<26> rd_sel<25> rs1_sel<25> rs2_sel<25> rd_sel<24> rs1_sel<24> rs2_sel<24> rd_sel<23>
+ rs1_sel<23> rs2_sel<23> rd_sel<22> rs1_sel<22> rs2_sel<22> rd_sel<21> rs1_sel<21> rs2_sel<21> rd_sel<20> rs1_sel<20> rs2_sel<20> rd_sel<19> rs1_sel<19> rs2_sel<19> rd_sel<18> rs1_sel<18> rs2_sel<18> rd_sel<17> rs1_sel<17> rs2_sel<17>
+ rd_sel<16> rs1_sel<16> rs2_sel<16> rd_sel<15> rs1_sel<15> rs2_sel<15> rd_sel<14> rs1_sel<14> rs2_sel<14> rd_sel<13> rs1_sel<13> rs2_sel<13> rd_sel<12> rs1_sel<12> rs2_sel<12> rd_sel<11> rs1_sel<11> rs2_sel<11> rd_sel<10> rs1_sel<10>
+ rs2_sel<10> rd_sel<9> rs1_sel<9> rs2_sel<9> rd_sel<8> rs1_sel<8> rs2_sel<8> rd_sel<7> rs1_sel<7> rs2_sel<7> rd_sel<6> rs1_sel<6> rs2_sel<6> rd_sel<5> rs1_sel<5> rs2_sel<5> rd_sel<4> rs1_sel<4> rs2_sel<4> rd_sel<3>
+ rs1_sel<3> rs2_sel<3> rd_sel<2> rs1_sel<2> rs2_sel<2> rd_sel<1> rs1_sel<1> rs2_sel<1> rs2_sel<0> rs1_sel<0> clk dmem_wdata<12> dmem_wdata<11> alu_mux_1_sel imem_addr<12> imem_addr<11> alu_inv_rs2 alu_mux_2_sel 324 shift_out<62>
+ alu_op<0> alu_op<1> shift_dir shift_out<55> shift_out<50> shift_out<65> shift_out<60> shift_out<51> shift_out<66> shift_out<46> shift_out<71> shift_out<42> 363 364 365 shift_out<23> shift_out<18> 368 shift_out<98> shift_out<144>
+ shift_out<139> 214 shift_out<61> shift_out<56> shift_amount<1> 372 shift_amount<2> shift_out<63> shift_out<58> shift_amount<3> 373 374 shift_amount<4> cmp_mux_sel 343 376 344 345 377 pc_mux_sel
+ rst 24 26
+ ICV_29 $T=0 0 0 0 $X=0 $Y=86200
X6 mem_mux_sel<0> dmem_rdata<14> dmem_rdata<13> dmem_rdata<7> 27 29 mem_mux_sel<1> mem_mux_sel<2> rd_mux_sel<0> imm<14> imm<13> dmem_addr<14> dmem_addr<13> rd_mux_sel<1> rd_mux_sel<2> rd_sel<31> rs1_sel<31> rs2_sel<31> rd_sel<30> rs1_sel<30>
+ rs2_sel<30> rd_sel<29> rs1_sel<29> rs2_sel<29> rd_sel<28> rs1_sel<28> rs2_sel<28> rd_sel<27> rs1_sel<27> rs2_sel<27> rd_sel<26> rs1_sel<26> rs2_sel<26> rd_sel<25> rs1_sel<25> rs2_sel<25> rd_sel<24> rs1_sel<24> rs2_sel<24> rd_sel<23>
+ rs1_sel<23> rs2_sel<23> rd_sel<22> rs1_sel<22> rs2_sel<22> rd_sel<21> rs1_sel<21> rs2_sel<21> rd_sel<20> rs1_sel<20> rs2_sel<20> rd_sel<19> rs1_sel<19> rs2_sel<19> rd_sel<18> rs1_sel<18> rs2_sel<18> rd_sel<17> rs1_sel<17> rs2_sel<17>
+ rd_sel<16> rs1_sel<16> rs2_sel<16> rd_sel<15> rs1_sel<15> rs2_sel<15> rd_sel<14> rs1_sel<14> rs2_sel<14> rd_sel<13> rs1_sel<13> rs2_sel<13> rd_sel<12> rs1_sel<12> rs2_sel<12> rd_sel<11> rs1_sel<11> rs2_sel<11> rd_sel<10> rs1_sel<10>
+ rs2_sel<10> rd_sel<9> rs1_sel<9> rs2_sel<9> rd_sel<8> rs1_sel<8> rs2_sel<8> rd_sel<7> rs1_sel<7> rs2_sel<7> rd_sel<6> rs1_sel<6> rs2_sel<6> rd_sel<5> rs1_sel<5> rs2_sel<5> rd_sel<4> rs1_sel<4> rs2_sel<4> rd_sel<3>
+ rs1_sel<3> rs2_sel<3> rd_sel<2> rs1_sel<2> rs2_sel<2> rd_sel<1> rs1_sel<1> rs2_sel<1> rs2_sel<0> rs1_sel<0> clk dmem_wdata<14> dmem_wdata<13> alu_mux_1_sel imem_addr<14> imem_addr<13> alu_inv_rs2 alu_mux_2_sel 354 386
+ shift_out<67> shift_out<72> alu_op<0> alu_op<1> shift_dir shift_out<65> shift_out<60> shift_out<75> shift_out<70> shift_out<61> shift_out<76> shift_out<56> shift_out<81> 395 396 397 398 shift_out<33> shift_out<28> 401
+ 402 shift_out<154> shift_out<149> 214 shift_out<71> shift_out<66> shift_amount<1> shift_amount<2> shift_out<73> shift_out<68> shift_amount<3> 405 406 shift_amount<4> cmp_mux_sel 375 408 376 377 409
+ pc_mux_sel rst 28 30
+ ICV_30 $T=0 0 0 0 $X=0 $Y=77000
X7 mem_mux_sel<0> dmem_rdata<16> dmem_rdata<15> dmem_rdata<7> 31 33 mem_mux_sel<1> mem_mux_sel<2> rd_mux_sel<0> imm<16> imm<15> dmem_addr<16> dmem_addr<15> shift_out<22> rd_mux_sel<1> rd_mux_sel<2> rd_sel<31> rs1_sel<31> rs2_sel<31> rd_sel<30>
+ rs1_sel<30> rs2_sel<30> rd_sel<29> rs1_sel<29> rs2_sel<29> rd_sel<28> rs1_sel<28> rs2_sel<28> rd_sel<27> rs1_sel<27> rs2_sel<27> rd_sel<26> rs1_sel<26> rs2_sel<26> rd_sel<25> rs1_sel<25> rs2_sel<25> rd_sel<24> rs1_sel<24> rs2_sel<24>
+ rd_sel<23> rs1_sel<23> rs2_sel<23> rd_sel<22> rs1_sel<22> rs2_sel<22> rd_sel<21> rs1_sel<21> rs2_sel<21> rd_sel<20> rs1_sel<20> rs2_sel<20> rd_sel<19> rs1_sel<19> rs2_sel<19> rd_sel<18> rs1_sel<18> rs2_sel<18> rd_sel<17> rs1_sel<17>
+ rs2_sel<17> rd_sel<16> rs1_sel<16> rs2_sel<16> rd_sel<15> rs1_sel<15> rs2_sel<15> rd_sel<14> rs1_sel<14> rs2_sel<14> rd_sel<13> rs1_sel<13> rs2_sel<13> rd_sel<12> rs1_sel<12> rs2_sel<12> rd_sel<11> rs1_sel<11> rs2_sel<11> rd_sel<10>
+ rs1_sel<10> rs2_sel<10> rd_sel<9> rs1_sel<9> rs2_sel<9> rd_sel<8> rs1_sel<8> rs2_sel<8> rd_sel<7> rs1_sel<7> rs2_sel<7> rd_sel<6> rs1_sel<6> rs2_sel<6> rd_sel<5> rs1_sel<5> rs2_sel<5> rd_sel<4> rs1_sel<4> rs2_sel<4>
+ rd_sel<3> rs1_sel<3> rs2_sel<3> rd_sel<2> rs1_sel<2> rs2_sel<2> rd_sel<1> rs1_sel<1> rs2_sel<1> rs2_sel<0> rs1_sel<0> clk dmem_wdata<16> dmem_wdata<15> alu_mux_1_sel imem_addr<16> imem_addr<15> alu_inv_rs2 alu_mux_2_sel 386
+ shift_out<82> shift_out<62> shift_out<77> alu_op<0> alu_op<1> shift_dir shift_out<75> shift_out<70> shift_out<85> shift_out<80> shift_out<71> shift_out<66> shift_out<91> shift_out<86> shift_out<57> 427 428 429 shift_out<38> shift_out<123>
+ 432 shift_out<4> shift_msb shift_out<159> 214 shift_out<81> shift_out<76> shift_amount<1> shift_amount<2> 437 438 shift_amount<3> shift_out<84> 440 shift_amount<4> cmp_mux_sel 407 442 408 409
+ 443 pc_mux_sel rst 32 34
+ ICV_31 $T=0 0 0 0 $X=0 $Y=67600
X8 mem_mux_sel<0> dmem_rdata<20> dmem_rdata<19> dmem_rdata<18> dmem_rdata<17> dmem_rdata<7> dmem_rdata<15> 35 37 39 41 mem_mux_sel<1> mem_mux_sel<2> rd_mux_sel<0> imm<20> imm<19> imm<18> imm<17> dmem_addr<20> dmem_addr<19>
+ dmem_addr<18> dmem_addr<17> shift_out<104> shift_out<99> shift_out<94> shift_out<89> rd_mux_sel<1> rd_mux_sel<2> rd_sel<31> rs1_sel<31> rs2_sel<31> rd_sel<30> rs1_sel<30> rs2_sel<30> rd_sel<29> rs1_sel<29> rs2_sel<29> rd_sel<28> rs1_sel<28> rs2_sel<28>
+ rd_sel<27> rs1_sel<27> rs2_sel<27> rd_sel<26> rs1_sel<26> rs2_sel<26> rd_sel<25> rs1_sel<25> rs2_sel<25> rd_sel<24> rs1_sel<24> rs2_sel<24> rd_sel<23> rs1_sel<23> rs2_sel<23> rd_sel<22> rs1_sel<22> rs2_sel<22> rd_sel<21> rs1_sel<21>
+ rs2_sel<21> rd_sel<20> rs1_sel<20> rs2_sel<20> rd_sel<19> rs1_sel<19> rs2_sel<19> rd_sel<18> rs1_sel<18> rs2_sel<18> rd_sel<17> rs1_sel<17> rs2_sel<17> rd_sel<16> rs1_sel<16> rs2_sel<16> rd_sel<15> rs1_sel<15> rs2_sel<15> rd_sel<14>
+ rs1_sel<14> rs2_sel<14> rd_sel<13> rs1_sel<13> rs2_sel<13> rd_sel<12> rs1_sel<12> rs2_sel<12> rd_sel<11> rs1_sel<11> rs2_sel<11> rd_sel<10> rs1_sel<10> rs2_sel<10> rd_sel<9> rs1_sel<9> rs2_sel<9> rd_sel<8> rs1_sel<8> rs2_sel<8>
+ rd_sel<7> rs1_sel<7> rs2_sel<7> rd_sel<6> rs1_sel<6> rs2_sel<6> rd_sel<5> rs1_sel<5> rs2_sel<5> rd_sel<4> rs1_sel<4> rs2_sel<4> rd_sel<3> rs1_sel<3> rs2_sel<3> rd_sel<2> rs1_sel<2> rs2_sel<2> rd_sel<1> rs1_sel<1>
+ rs2_sel<1> rs2_sel<0> rs1_sel<0> clk dmem_wdata<20> dmem_wdata<19> dmem_wdata<18> dmem_wdata<17> alu_mux_1_sel imem_addr<20> imem_addr<19> imem_addr<18> imem_addr<17> alu_inv_rs2 alu_mux_2_sel 418 458 shift_out<82> shift_out<87> shift_out<92>
+ shift_out<72> shift_out<97> shift_out<77> alu_op<0> alu_op<1> shift_dir shift_out<95> shift_out<90> shift_out<85> shift_out<80> shift_out<105> shift_out<100> shift_out<91> shift_out<106> shift_out<86> shift_out<81> shift_out<96> shift_out<76> shift_out<111> shift_out<101>
+ shift_out<67> 474 475 476 477 478 479 480 481 shift_out<143> shift_out<138> shift_out<133> shift_out<128> shift_out<24> shift_out<19> shift_out<14> shift_out<9> shift_msb 214 shift_amount<1>
+ shift_out<102> shift_amount<2> 491 492 493 494 shift_amount<3> 495 496 497 498 shift_amount<4> cmp_mux_sel 499 441 500 442 443 501 pc_mux_sel
+ rst 36 38 40 42
+ ICV_36 $T=0 0 0 0 $X=0 $Y=50930
X9 mem_mux_sel<0> dmem_rdata<22> dmem_rdata<21> dmem_rdata<7> dmem_rdata<15> 43 45 mem_mux_sel<1> mem_mux_sel<2> rd_mux_sel<0> imm<22> imm<21> dmem_addr<22> dmem_addr<21> shift_out<114> shift_out<109> rd_mux_sel<1> rd_mux_sel<2> rd_sel<31> rs1_sel<31>
+ rs2_sel<31> rd_sel<30> rs1_sel<30> rs2_sel<30> rd_sel<29> rs1_sel<29> rs2_sel<29> rd_sel<28> rs1_sel<28> rs2_sel<28> rd_sel<27> rs1_sel<27> rs2_sel<27> rd_sel<26> rs1_sel<26> rs2_sel<26> rd_sel<25> rs1_sel<25> rs2_sel<25> rd_sel<24>
+ rs1_sel<24> rs2_sel<24> rd_sel<23> rs1_sel<23> rs2_sel<23> rd_sel<22> rs1_sel<22> rs2_sel<22> rd_sel<21> rs1_sel<21> rs2_sel<21> rd_sel<20> rs1_sel<20> rs2_sel<20> rd_sel<19> rs1_sel<19> rs2_sel<19> rd_sel<18> rs1_sel<18> rs2_sel<18>
+ rd_sel<17> rs1_sel<17> rs2_sel<17> rd_sel<16> rs1_sel<16> rs2_sel<16> rd_sel<15> rs1_sel<15> rs2_sel<15> rd_sel<14> rs1_sel<14> rs2_sel<14> rd_sel<13> rs1_sel<13> rs2_sel<13> rd_sel<12> rs1_sel<12> rs2_sel<12> rd_sel<11> rs1_sel<11>
+ rs2_sel<11> rd_sel<10> rs1_sel<10> rs2_sel<10> rd_sel<9> rs1_sel<9> rs2_sel<9> rd_sel<8> rs1_sel<8> rs2_sel<8> rd_sel<7> rs1_sel<7> rs2_sel<7> rd_sel<6> rs1_sel<6> rs2_sel<6> rd_sel<5> rs1_sel<5> rs2_sel<5> rd_sel<4>
+ rs1_sel<4> rs2_sel<4> rd_sel<3> rs1_sel<3> rs2_sel<3> rd_sel<2> rs1_sel<2> rs2_sel<2> rd_sel<1> rs1_sel<1> rs2_sel<1> rs2_sel<0> rs1_sel<0> clk dmem_wdata<22> dmem_wdata<21> alu_mux_1_sel imem_addr<22> imem_addr<21> alu_inv_rs2
+ alu_mux_2_sel 512 shift_out<107> shift_out<87> shift_out<92> alu_op<0> alu_op<1> shift_dir shift_out<105> shift_out<100> shift_out<115> shift_out<110> shift_out<101> shift_out<116> shift_out<96> shift_out<121> 520 521 522 523
+ shift_out<153> shift_out<148> shift_out<34> shift_out<29> shift_msb 214 shift_out<111> shift_out<106> shift_amount<1> shift_out<112> shift_amount<2> 529 530 shift_amount<3> 531 532 shift_amount<4> cmp_mux_sel 66 67
+ 500 501 534 pc_mux_sel rst 44 46
+ ICV_37 $T=0 0 0 0 $X=0 $Y=41600
X10 mem_mux_sel<0> dmem_rdata<24> dmem_rdata<23> dmem_rdata<7> dmem_rdata<15> 47 49 mem_mux_sel<1> mem_mux_sel<2> rd_mux_sel<0> imm<24> imm<23> dmem_addr<24> dmem_addr<23> rd_mux_sel<1> rd_mux_sel<2> rd_sel<31> rs1_sel<31> rs2_sel<31> rd_sel<30>
+ rs1_sel<30> rs2_sel<30> rd_sel<29> rs1_sel<29> rs2_sel<29> rd_sel<28> rs1_sel<28> rs2_sel<28> rd_sel<27> rs1_sel<27> rs2_sel<27> rd_sel<26> rs1_sel<26> rs2_sel<26> rd_sel<25> rs1_sel<25> rs2_sel<25> rd_sel<24> rs1_sel<24> rs2_sel<24>
+ rd_sel<23> rs1_sel<23> rs2_sel<23> rd_sel<22> rs1_sel<22> rs2_sel<22> rd_sel<21> rs1_sel<21> rs2_sel<21> rd_sel<20> rs1_sel<20> rs2_sel<20> rd_sel<19> rs1_sel<19> rs2_sel<19> rd_sel<18> rs1_sel<18> rs2_sel<18> rd_sel<17> rs1_sel<17>
+ rs2_sel<17> rd_sel<16> rs1_sel<16> rs2_sel<16> rd_sel<15> rs1_sel<15> rs2_sel<15> rd_sel<14> rs1_sel<14> rs2_sel<14> rd_sel<13> rs1_sel<13> rs2_sel<13> rd_sel<12> rs1_sel<12> rs2_sel<12> rd_sel<11> rs1_sel<11> rs2_sel<11> rd_sel<10>
+ rs1_sel<10> rs2_sel<10> rd_sel<9> rs1_sel<9> rs2_sel<9> rd_sel<8> rs1_sel<8> rs2_sel<8> rd_sel<7> rs1_sel<7> rs2_sel<7> rd_sel<6> rs1_sel<6> rs2_sel<6> rd_sel<5> rs1_sel<5> rs2_sel<5> rd_sel<4> rs1_sel<4> rs2_sel<4>
+ rd_sel<3> rs1_sel<3> rs2_sel<3> rd_sel<2> rs1_sel<2> rs2_sel<2> rd_sel<1> rs1_sel<1> rs2_sel<1> rs2_sel<0> rs1_sel<0> clk dmem_wdata<24> dmem_wdata<23> alu_mux_1_sel imem_addr<24> imem_addr<23> alu_inv_rs2 alu_mux_2_sel 512
+ 543 shift_out<102> shift_out<117> shift_out<97> alu_op<0> alu_op<1> shift_dir shift_out<115> shift_out<110> shift_out<125> shift_out<120> shift_out<111> shift_out<126> shift_out<106> shift_out<131> shift_out<142> 552 shift_out<83> shift_out<78> shift_msb
+ shift_out<158> shift_out<44> shift_out<39> 214 shift_out<121> shift_out<116> shift_amount<1> shift_out<122> shift_amount<2> 559 560 shift_amount<3> 561 562 shift_amount<4> cmp_mux_sel 563 533 68 67
+ 534 564 pc_mux_sel rst 48 50
+ ICV_38 $T=0 0 0 0 $X=0 $Y=32400
X11 mem_mux_sel<0> dmem_rdata<26> dmem_rdata<25> dmem_rdata<7> dmem_rdata<15> 51 53 mem_mux_sel<1> mem_mux_sel<2> rd_mux_sel<0> imm<26> imm<25> dmem_addr<26> dmem_addr<25> rd_mux_sel<1> rd_mux_sel<2> rd_sel<31> rs1_sel<31> rs2_sel<31> rd_sel<30>
+ rs1_sel<30> rs2_sel<30> rd_sel<29> rs1_sel<29> rs2_sel<29> rd_sel<28> rs1_sel<28> rs2_sel<28> rd_sel<27> rs1_sel<27> rs2_sel<27> rd_sel<26> rs1_sel<26> rs2_sel<26> rd_sel<25> rs1_sel<25> rs2_sel<25> rd_sel<24> rs1_sel<24> rs2_sel<24>
+ rd_sel<23> rs1_sel<23> rs2_sel<23> rd_sel<22> rs1_sel<22> rs2_sel<22> rd_sel<21> rs1_sel<21> rs2_sel<21> rd_sel<20> rs1_sel<20> rs2_sel<20> rd_sel<19> rs1_sel<19> rs2_sel<19> rd_sel<18> rs1_sel<18> rs2_sel<18> rd_sel<17> rs1_sel<17>
+ rs2_sel<17> rd_sel<16> rs1_sel<16> rs2_sel<16> rd_sel<15> rs1_sel<15> rs2_sel<15> rd_sel<14> rs1_sel<14> rs2_sel<14> rd_sel<13> rs1_sel<13> rs2_sel<13> rd_sel<12> rs1_sel<12> rs2_sel<12> rd_sel<11> rs1_sel<11> rs2_sel<11> rd_sel<10>
+ rs1_sel<10> rs2_sel<10> rd_sel<9> rs1_sel<9> rs2_sel<9> rd_sel<8> rs1_sel<8> rs2_sel<8> rd_sel<7> rs1_sel<7> rs2_sel<7> rd_sel<6> rs1_sel<6> rs2_sel<6> rd_sel<5> rs1_sel<5> rs2_sel<5> rd_sel<4> rs1_sel<4> rs2_sel<4>
+ rd_sel<3> rs1_sel<3> rs2_sel<3> rd_sel<2> rs1_sel<2> rs2_sel<2> rd_sel<1> rs1_sel<1> rs2_sel<1> rs2_sel<0> rs1_sel<0> clk dmem_wdata<26> dmem_wdata<25> alu_mux_1_sel imem_addr<26> imem_addr<25> alu_inv_rs2 alu_mux_2_sel 573
+ shift_out<127> shift_out<107> shift_out<112> alu_op<0> alu_op<1> shift_dir shift_out<125> shift_out<120> shift_out<135> shift_out<130> shift_out<121> shift_out<136> shift_out<116> shift_out<141> shift_out<152> shift_out<147> shift_out<93> shift_out<88> shift_msb shift_out<54>
+ shift_out<49> 214 shift_out<131> shift_out<126> shift_amount<1> shift_out<132> shift_amount<2> 588 589 shift_amount<3> 590 591 shift_amount<4> cmp_mux_sel 592 593 68 564 594 pc_mux_sel
+ rst 52 54
+ ICV_39 $T=0 0 0 0 $X=0 $Y=23150
X12 mem_mux_sel<0> dmem_rdata<28> dmem_rdata<27> dmem_rdata<7> dmem_rdata<15> 55 57 mem_mux_sel<1> mem_mux_sel<2> rd_mux_sel<0> imm<28> imm<27> dmem_addr<28> dmem_addr<27> rd_mux_sel<1> rd_mux_sel<2> rd_sel<31> rs1_sel<31> rs2_sel<31> rd_sel<30>
+ rs1_sel<30> rs2_sel<30> rd_sel<29> rs1_sel<29> rs2_sel<29> rd_sel<28> rs1_sel<28> rs2_sel<28> rd_sel<27> rs1_sel<27> rs2_sel<27> rd_sel<26> rs1_sel<26> rs2_sel<26> rd_sel<25> rs1_sel<25> rs2_sel<25> rd_sel<24> rs1_sel<24> rs2_sel<24>
+ rd_sel<23> rs1_sel<23> rs2_sel<23> rd_sel<22> rs1_sel<22> rs2_sel<22> rd_sel<21> rs1_sel<21> rs2_sel<21> rd_sel<20> rs1_sel<20> rs2_sel<20> rd_sel<19> rs1_sel<19> rs2_sel<19> rd_sel<18> rs1_sel<18> rs2_sel<18> rd_sel<17> rs1_sel<17>
+ rs2_sel<17> rd_sel<16> rs1_sel<16> rs2_sel<16> rd_sel<15> rs1_sel<15> rs2_sel<15> rd_sel<14> rs1_sel<14> rs2_sel<14> rd_sel<13> rs1_sel<13> rs2_sel<13> rd_sel<12> rs1_sel<12> rs2_sel<12> rd_sel<11> rs1_sel<11> rs2_sel<11> rd_sel<10>
+ rs1_sel<10> rs2_sel<10> rd_sel<9> rs1_sel<9> rs2_sel<9> rd_sel<8> rs1_sel<8> rs2_sel<8> rd_sel<7> rs1_sel<7> rs2_sel<7> rd_sel<6> rs1_sel<6> rs2_sel<6> rd_sel<5> rs1_sel<5> rs2_sel<5> rd_sel<4> rs1_sel<4> rs2_sel<4>
+ rd_sel<3> rs1_sel<3> rs2_sel<3> rd_sel<2> rs1_sel<2> rs2_sel<2> rd_sel<1> rs1_sel<1> rs2_sel<1> rs2_sel<0> rs1_sel<0> clk dmem_wdata<28> dmem_wdata<27> alu_mux_1_sel imem_addr<28> imem_addr<27> alu_inv_rs2 alu_mux_2_sel 573
+ 603 shift_out<122> shift_out<137> shift_out<117> alu_op<0> alu_op<1> shift_dir shift_out<135> shift_out<130> shift_out<145> shift_out<140> shift_out<131> shift_out<146> shift_out<126> shift_out<151> shift_msb shift_out<157> shift_out<103> shift_out98> shift_out<64>
+ shift_out<59> 214 shift_out<141> shift_out<136> shift_amount<1> 616 shift_amount<2> 617 618 shift_amount<3> 619 620 shift_amount<4> cmp_mux_sel 69 70 593 594 622 pc_mux_sel
+ rst 56 58
+ ICV_40 $T=0 0 0 0 $X=0 $Y=13800
X13 mem_mux_sel<0> dmem_rdata<31> dmem_rdata<30> dmem_rdata<29> dmem_rdata<7> dmem_rdata<15> vss! 61 63 mem_mux_sel<1> mem_mux_sel<2> rd_mux_sel<0> imm<31> imm<30> imm<29> dmem_addr<31> dmem_addr<30> dmem_addr<29> rd_mux_sel<1> rd_mux_sel<2>
+ rd_sel<31> rs1_sel<31> rs2_sel<31> rd_sel<30> rs1_sel<30> rs2_sel<30> rd_sel<29> rs1_sel<29> rs2_sel<29> rd_sel<28> rs1_sel<28> rs2_sel<28> rd_sel<27> rs1_sel<27> rs2_sel<27> rd_sel<26> rs1_sel<26> rs2_sel<26> rd_sel<25> rs1_sel<25>
+ rs2_sel<25> rd_sel<24> rs1_sel<24> rs2_sel<24> rd_sel<23> rs1_sel<23> rs2_sel<23> rd_sel<22> rs1_sel<22> rs2_sel<22> rd_sel<21> rs1_sel<21> rs2_sel<21> rd_sel<20> rs1_sel<20> rs2_sel<20> rd_sel<19> rs1_sel<19> rs2_sel<19> rd_sel<18>
+ rs1_sel<18> rs2_sel<18> rd_sel<17> rs1_sel<17> rs2_sel<17> rd_sel<16> rs1_sel<16> rs2_sel<16> rd_sel<15> rs1_sel<15> rs2_sel<15> rd_sel<14> rs1_sel<14> rs2_sel<14> rd_sel<13> rs1_sel<13> rs2_sel<13> rd_sel<12> rs1_sel<12> rs2_sel<12>
+ rd_sel<11> rs1_sel<11> rs2_sel<11> rd_sel<10> rs1_sel<10> rs2_sel<10> rd_sel<9> rs1_sel<9> rs2_sel<9> rd_sel<8> rs1_sel<8> rs2_sel<8> rd_sel<7> rs1_sel<7> rs2_sel<7> rd_sel<6> rs1_sel<6> rs2_sel<6> rd_sel<5> rs1_sel<5>
+ rs2_sel<5> rd_sel<4> rs1_sel<4> rs2_sel<4> rd_sel<3> rs1_sel<3> rs2_sel<3> rd_sel<2> rs1_sel<2> rs2_sel<2> rd_sel<1> rs1_sel<1> rs2_sel<1> rs2_sel<0> rs1_sel<0> clk cmp_a_31 dmem_wdata<31> dmem_wdata<30> dmem_wdata<29>
+ alu_mux_1_sel imem_addr<31> imem_addr<30> imem_addr<29> alu_inv_rs2 alu_mux_2_sel shift_out<127> shift_out<132> shift_out<137> alu_op<0> alu_op<1> shift_dir shift_out<150> shift_out<145> shift_out<140> shift_msb shift_out<155> shift_out<146> shift_out<141> shift_out<136>
+ shift_out<156> shift_out<118> shift_out<113> shift_out<108> shift_out<79> shift_out<74> shift_out<69> 214 646 shift_out<151> shift_amount<1> 647 648 649 shift_amount<2> 650 651 652 shift_amount<3> 653
+ 654 655 shift_amount<4> cmp_mux_sel cmp_b_31 vdd! 621 70 622 pc_mux_sel rst 62 64
+ ICV_41 $T=0 0 0 0 $X=0 $Y=0
*.CALIBRE WARNING SHORT Short circuit(s) detected by extraction in this cell. See extraction report for details.
*.CALIBRE WARNING OPEN Open circuit(s) detected by extraction in this cell. See extraction report for details.
.ENDS
***************************************
